// 1 2 1 2 1 2 2 1 2 1 1 1 2 2 2 1 2 2 1 2 2 1 2 2 2 2 2 2 2 2 2 2 

module main(x,y,o);
input [15:0] x,y;
output [31:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_1_0,x[1],y[0]);
and and17(ip_1_1,x[1],y[1]);
and and18(ip_1_2,x[1],y[2]);
and and19(ip_1_3,x[1],y[3]);
and and20(ip_1_4,x[1],y[4]);
and and21(ip_1_5,x[1],y[5]);
and and22(ip_1_6,x[1],y[6]);
and and23(ip_1_7,x[1],y[7]);
and and24(ip_1_8,x[1],y[8]);
and and25(ip_1_9,x[1],y[9]);
and and26(ip_1_10,x[1],y[10]);
and and27(ip_1_11,x[1],y[11]);
and and28(ip_1_12,x[1],y[12]);
and and29(ip_1_13,x[1],y[13]);
and and30(ip_1_14,x[1],y[14]);
and and31(ip_1_15,x[1],y[15]);
and and32(ip_2_0,x[2],y[0]);
and and33(ip_2_1,x[2],y[1]);
and and34(ip_2_2,x[2],y[2]);
and and35(ip_2_3,x[2],y[3]);
and and36(ip_2_4,x[2],y[4]);
and and37(ip_2_5,x[2],y[5]);
and and38(ip_2_6,x[2],y[6]);
and and39(ip_2_7,x[2],y[7]);
and and40(ip_2_8,x[2],y[8]);
and and41(ip_2_9,x[2],y[9]);
and and42(ip_2_10,x[2],y[10]);
and and43(ip_2_11,x[2],y[11]);
and and44(ip_2_12,x[2],y[12]);
and and45(ip_2_13,x[2],y[13]);
and and46(ip_2_14,x[2],y[14]);
and and47(ip_2_15,x[2],y[15]);
and and48(ip_3_0,x[3],y[0]);
and and49(ip_3_1,x[3],y[1]);
and and50(ip_3_2,x[3],y[2]);
and and51(ip_3_3,x[3],y[3]);
and and52(ip_3_4,x[3],y[4]);
and and53(ip_3_5,x[3],y[5]);
and and54(ip_3_6,x[3],y[6]);
and and55(ip_3_7,x[3],y[7]);
and and56(ip_3_8,x[3],y[8]);
and and57(ip_3_9,x[3],y[9]);
and and58(ip_3_10,x[3],y[10]);
and and59(ip_3_11,x[3],y[11]);
and and60(ip_3_12,x[3],y[12]);
and and61(ip_3_13,x[3],y[13]);
and and62(ip_3_14,x[3],y[14]);
and and63(ip_3_15,x[3],y[15]);
and and64(ip_4_0,x[4],y[0]);
and and65(ip_4_1,x[4],y[1]);
and and66(ip_4_2,x[4],y[2]);
and and67(ip_4_3,x[4],y[3]);
and and68(ip_4_4,x[4],y[4]);
and and69(ip_4_5,x[4],y[5]);
and and70(ip_4_6,x[4],y[6]);
and and71(ip_4_7,x[4],y[7]);
and and72(ip_4_8,x[4],y[8]);
and and73(ip_4_9,x[4],y[9]);
and and74(ip_4_10,x[4],y[10]);
and and75(ip_4_11,x[4],y[11]);
and and76(ip_4_12,x[4],y[12]);
and and77(ip_4_13,x[4],y[13]);
and and78(ip_4_14,x[4],y[14]);
and and79(ip_4_15,x[4],y[15]);
and and80(ip_5_0,x[5],y[0]);
and and81(ip_5_1,x[5],y[1]);
and and82(ip_5_2,x[5],y[2]);
and and83(ip_5_3,x[5],y[3]);
and and84(ip_5_4,x[5],y[4]);
and and85(ip_5_5,x[5],y[5]);
and and86(ip_5_6,x[5],y[6]);
and and87(ip_5_7,x[5],y[7]);
and and88(ip_5_8,x[5],y[8]);
and and89(ip_5_9,x[5],y[9]);
and and90(ip_5_10,x[5],y[10]);
and and91(ip_5_11,x[5],y[11]);
and and92(ip_5_12,x[5],y[12]);
and and93(ip_5_13,x[5],y[13]);
and and94(ip_5_14,x[5],y[14]);
and and95(ip_5_15,x[5],y[15]);
and and96(ip_6_0,x[6],y[0]);
and and97(ip_6_1,x[6],y[1]);
and and98(ip_6_2,x[6],y[2]);
and and99(ip_6_3,x[6],y[3]);
and and100(ip_6_4,x[6],y[4]);
and and101(ip_6_5,x[6],y[5]);
and and102(ip_6_6,x[6],y[6]);
and and103(ip_6_7,x[6],y[7]);
and and104(ip_6_8,x[6],y[8]);
and and105(ip_6_9,x[6],y[9]);
and and106(ip_6_10,x[6],y[10]);
and and107(ip_6_11,x[6],y[11]);
and and108(ip_6_12,x[6],y[12]);
and and109(ip_6_13,x[6],y[13]);
and and110(ip_6_14,x[6],y[14]);
and and111(ip_6_15,x[6],y[15]);
and and112(ip_7_0,x[7],y[0]);
and and113(ip_7_1,x[7],y[1]);
and and114(ip_7_2,x[7],y[2]);
and and115(ip_7_3,x[7],y[3]);
and and116(ip_7_4,x[7],y[4]);
and and117(ip_7_5,x[7],y[5]);
and and118(ip_7_6,x[7],y[6]);
and and119(ip_7_7,x[7],y[7]);
and and120(ip_7_8,x[7],y[8]);
and and121(ip_7_9,x[7],y[9]);
and and122(ip_7_10,x[7],y[10]);
and and123(ip_7_11,x[7],y[11]);
and and124(ip_7_12,x[7],y[12]);
and and125(ip_7_13,x[7],y[13]);
and and126(ip_7_14,x[7],y[14]);
and and127(ip_7_15,x[7],y[15]);
and and128(ip_8_0,x[8],y[0]);
and and129(ip_8_1,x[8],y[1]);
and and130(ip_8_2,x[8],y[2]);
and and131(ip_8_3,x[8],y[3]);
and and132(ip_8_4,x[8],y[4]);
and and133(ip_8_5,x[8],y[5]);
and and134(ip_8_6,x[8],y[6]);
and and135(ip_8_7,x[8],y[7]);
and and136(ip_8_8,x[8],y[8]);
and and137(ip_8_9,x[8],y[9]);
and and138(ip_8_10,x[8],y[10]);
and and139(ip_8_11,x[8],y[11]);
and and140(ip_8_12,x[8],y[12]);
and and141(ip_8_13,x[8],y[13]);
and and142(ip_8_14,x[8],y[14]);
and and143(ip_8_15,x[8],y[15]);
and and144(ip_9_0,x[9],y[0]);
and and145(ip_9_1,x[9],y[1]);
and and146(ip_9_2,x[9],y[2]);
and and147(ip_9_3,x[9],y[3]);
and and148(ip_9_4,x[9],y[4]);
and and149(ip_9_5,x[9],y[5]);
and and150(ip_9_6,x[9],y[6]);
and and151(ip_9_7,x[9],y[7]);
and and152(ip_9_8,x[9],y[8]);
and and153(ip_9_9,x[9],y[9]);
and and154(ip_9_10,x[9],y[10]);
and and155(ip_9_11,x[9],y[11]);
and and156(ip_9_12,x[9],y[12]);
and and157(ip_9_13,x[9],y[13]);
and and158(ip_9_14,x[9],y[14]);
and and159(ip_9_15,x[9],y[15]);
and and160(ip_10_0,x[10],y[0]);
and and161(ip_10_1,x[10],y[1]);
and and162(ip_10_2,x[10],y[2]);
and and163(ip_10_3,x[10],y[3]);
and and164(ip_10_4,x[10],y[4]);
and and165(ip_10_5,x[10],y[5]);
and and166(ip_10_6,x[10],y[6]);
and and167(ip_10_7,x[10],y[7]);
and and168(ip_10_8,x[10],y[8]);
and and169(ip_10_9,x[10],y[9]);
and and170(ip_10_10,x[10],y[10]);
and and171(ip_10_11,x[10],y[11]);
and and172(ip_10_12,x[10],y[12]);
and and173(ip_10_13,x[10],y[13]);
and and174(ip_10_14,x[10],y[14]);
and and175(ip_10_15,x[10],y[15]);
and and176(ip_11_0,x[11],y[0]);
and and177(ip_11_1,x[11],y[1]);
and and178(ip_11_2,x[11],y[2]);
and and179(ip_11_3,x[11],y[3]);
and and180(ip_11_4,x[11],y[4]);
and and181(ip_11_5,x[11],y[5]);
and and182(ip_11_6,x[11],y[6]);
and and183(ip_11_7,x[11],y[7]);
and and184(ip_11_8,x[11],y[8]);
and and185(ip_11_9,x[11],y[9]);
and and186(ip_11_10,x[11],y[10]);
and and187(ip_11_11,x[11],y[11]);
and and188(ip_11_12,x[11],y[12]);
and and189(ip_11_13,x[11],y[13]);
and and190(ip_11_14,x[11],y[14]);
and and191(ip_11_15,x[11],y[15]);
and and192(ip_12_0,x[12],y[0]);
and and193(ip_12_1,x[12],y[1]);
and and194(ip_12_2,x[12],y[2]);
and and195(ip_12_3,x[12],y[3]);
and and196(ip_12_4,x[12],y[4]);
and and197(ip_12_5,x[12],y[5]);
and and198(ip_12_6,x[12],y[6]);
and and199(ip_12_7,x[12],y[7]);
and and200(ip_12_8,x[12],y[8]);
and and201(ip_12_9,x[12],y[9]);
and and202(ip_12_10,x[12],y[10]);
and and203(ip_12_11,x[12],y[11]);
and and204(ip_12_12,x[12],y[12]);
and and205(ip_12_13,x[12],y[13]);
and and206(ip_12_14,x[12],y[14]);
and and207(ip_12_15,x[12],y[15]);
and and208(ip_13_0,x[13],y[0]);
and and209(ip_13_1,x[13],y[1]);
and and210(ip_13_2,x[13],y[2]);
and and211(ip_13_3,x[13],y[3]);
and and212(ip_13_4,x[13],y[4]);
and and213(ip_13_5,x[13],y[5]);
and and214(ip_13_6,x[13],y[6]);
and and215(ip_13_7,x[13],y[7]);
and and216(ip_13_8,x[13],y[8]);
and and217(ip_13_9,x[13],y[9]);
and and218(ip_13_10,x[13],y[10]);
and and219(ip_13_11,x[13],y[11]);
and and220(ip_13_12,x[13],y[12]);
and and221(ip_13_13,x[13],y[13]);
and and222(ip_13_14,x[13],y[14]);
and and223(ip_13_15,x[13],y[15]);
and and224(ip_14_0,x[14],y[0]);
and and225(ip_14_1,x[14],y[1]);
and and226(ip_14_2,x[14],y[2]);
and and227(ip_14_3,x[14],y[3]);
and and228(ip_14_4,x[14],y[4]);
and and229(ip_14_5,x[14],y[5]);
and and230(ip_14_6,x[14],y[6]);
and and231(ip_14_7,x[14],y[7]);
and and232(ip_14_8,x[14],y[8]);
and and233(ip_14_9,x[14],y[9]);
and and234(ip_14_10,x[14],y[10]);
and and235(ip_14_11,x[14],y[11]);
and and236(ip_14_12,x[14],y[12]);
and and237(ip_14_13,x[14],y[13]);
and and238(ip_14_14,x[14],y[14]);
and and239(ip_14_15,x[14],y[15]);
and and240(ip_15_0,x[15],y[0]);
and and241(ip_15_1,x[15],y[1]);
and and242(ip_15_2,x[15],y[2]);
and and243(ip_15_3,x[15],y[3]);
and and244(ip_15_4,x[15],y[4]);
and and245(ip_15_5,x[15],y[5]);
and and246(ip_15_6,x[15],y[6]);
and and247(ip_15_7,x[15],y[7]);
and and248(ip_15_8,x[15],y[8]);
and and249(ip_15_9,x[15],y[9]);
and and250(ip_15_10,x[15],y[10]);
and and251(ip_15_11,x[15],y[11]);
and and252(ip_15_12,x[15],y[12]);
and and253(ip_15_13,x[15],y[13]);
and and254(ip_15_14,x[15],y[14]);
and and255(ip_15_15,x[15],y[15]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
HA ha0(ip_3_0,p3,p4,p5);
FA fa2(ip_0_4,ip_1_3,ip_2_2,p6,p7);
HA ha1(ip_3_1,ip_4_0,p8,p9);
HA ha2(p9,p7,p10,p11);
FA fa3(p11,p2,p4,p12,p13);
FA fa4(ip_0_5,ip_1_4,ip_2_3,p14,p15);
HA ha3(ip_3_2,ip_4_1,p16,p17);
HA ha4(ip_5_0,p17,p18,p19);
HA ha5(p8,p15,p20,p21);
FA fa5(p19,p10,p21,p22,p23);
HA ha6(p6,p23,p24,p25);
FA fa6(ip_0_6,ip_1_5,ip_2_4,p26,p27);
FA fa7(ip_3_3,ip_4_2,ip_5_1,p28,p29);
FA fa8(ip_6_0,p16,p18,p30,p31);
HA ha7(p27,p29,p32,p33);
FA fa9(p14,p20,p31,p34,p35);
FA fa10(p33,p35,p22,p36,p37);
HA ha8(ip_0_7,ip_1_6,p38,p39);
HA ha9(ip_2_5,ip_3_4,p40,p41);
FA fa11(ip_4_3,ip_5_2,ip_6_1,p42,p43);
FA fa12(ip_7_0,p39,p41,p44,p45);
FA fa13(p43,p26,p28,p46,p47);
HA ha10(p32,p45,p48,p49);
FA fa14(p30,p49,p47,p50,p51);
FA fa15(p34,p51,p36,p52,p53);
FA fa16(ip_0_8,ip_1_7,ip_2_6,p54,p55);
FA fa17(ip_3_5,ip_4_4,ip_5_3,p56,p57);
HA ha11(ip_6_2,ip_7_1,p58,p59);
FA fa18(ip_8_0,p38,p40,p60,p61);
HA ha12(p59,p55,p62,p63);
FA fa19(p57,p42,p61,p64,p65);
FA fa20(p63,p44,p48,p66,p67);
FA fa21(p65,p46,p67,p68,p69);
HA ha13(p50,p69,p70,p71);
FA fa22(ip_0_9,ip_1_8,ip_2_7,p72,p73);
FA fa23(ip_3_6,ip_4_5,ip_5_4,p74,p75);
HA ha14(ip_6_3,ip_7_2,p76,p77);
HA ha15(ip_8_1,ip_9_0,p78,p79);
FA fa24(p58,p77,p79,p80,p81);
FA fa25(p73,p75,p54,p82,p83);
HA ha16(p56,p62,p84,p85);
HA ha17(p81,p60,p86,p87);
FA fa26(p83,p85,p87,p88,p89);
FA fa27(p64,p89,p66,p90,p91);
FA fa28(p91,p68,p70,p92,p93);
FA fa29(ip_0_10,ip_1_9,ip_2_8,p94,p95);
FA fa30(ip_3_7,ip_4_6,ip_5_5,p96,p97);
FA fa31(ip_6_4,ip_7_3,ip_8_2,p98,p99);
FA fa32(ip_9_1,ip_10_0,p76,p100,p101);
FA fa33(p78,p101,p95,p102,p103);
HA ha18(p97,p99,p104,p105);
FA fa34(p105,p72,p74,p106,p107);
FA fa35(p103,p80,p84,p108,p109);
FA fa36(p107,p82,p86,p110,p111);
HA ha19(p109,p111,p112,p113);
HA ha20(p88,p113,p114,p115);
FA fa37(p115,p90,p92,p116,p117);
HA ha21(ip_0_11,ip_1_10,p118,p119);
FA fa38(ip_2_9,ip_3_8,ip_4_7,p120,p121);
FA fa39(ip_5_6,ip_6_5,ip_7_4,p122,p123);
HA ha22(ip_8_3,ip_9_2,p124,p125);
HA ha23(ip_10_1,ip_11_0,p126,p127);
HA ha24(p119,p125,p128,p129);
FA fa40(p127,p121,p123,p130,p131);
HA ha25(p129,p100,p132,p133);
HA ha26(p104,p94,p134,p135);
FA fa41(p96,p98,p131,p136,p137);
HA ha27(p133,p135,p138,p139);
HA ha28(p102,p137,p140,p141);
HA ha29(p139,p106,p142,p143);
FA fa42(p141,p108,p143,p144,p145);
FA fa43(p110,p112,p114,p146,p147);
FA fa44(p145,p147,p116,p148,p149);
FA fa45(ip_0_12,ip_1_11,ip_2_10,p150,p151);
FA fa46(ip_3_9,ip_4_8,ip_5_7,p152,p153);
FA fa47(ip_6_6,ip_7_5,ip_8_4,p154,p155);
FA fa48(ip_9_3,ip_10_2,ip_11_1,p156,p157);
FA fa49(ip_12_0,p118,p124,p158,p159);
FA fa50(p126,p128,p151,p160,p161);
HA ha30(p153,p155,p162,p163);
FA fa51(p157,p120,p122,p164,p165);
FA fa52(p159,p163,p132,p166,p167);
FA fa53(p134,p161,p130,p168,p169);
FA fa54(p138,p165,p167,p170,p171);
FA fa55(p136,p140,p169,p172,p173);
HA ha31(p142,p171,p174,p175);
HA ha32(p173,p175,p176,p177);
FA fa56(p177,p144,p146,p178,p179);
HA ha33(ip_0_13,ip_1_12,p180,p181);
FA fa57(ip_2_11,ip_3_10,ip_4_9,p182,p183);
HA ha34(ip_5_8,ip_6_7,p184,p185);
FA fa58(ip_7_6,ip_8_5,ip_9_4,p186,p187);
FA fa59(ip_10_3,ip_11_2,ip_12_1,p188,p189);
HA ha35(ip_13_0,p181,p190,p191);
FA fa60(p185,p183,p187,p192,p193);
HA ha36(p189,p191,p194,p195);
HA ha37(p150,p152,p196,p197);
HA ha38(p154,p156,p198,p199);
FA fa61(p162,p195,p158,p200,p201);
FA fa62(p193,p197,p199,p202,p203);
FA fa63(p160,p201,p164,p204,p205);
FA fa64(p166,p203,p168,p206,p207);
FA fa65(p205,p170,p174,p208,p209);
FA fa66(p207,p172,p176,p210,p211);
HA ha39(p209,p211,p212,p213);
HA ha40(ip_0_14,ip_1_13,p214,p215);
FA fa67(ip_2_12,ip_3_11,ip_4_10,p216,p217);
FA fa68(ip_5_9,ip_6_8,ip_7_7,p218,p219);
HA ha41(ip_8_6,ip_9_5,p220,p221);
HA ha42(ip_10_4,ip_11_3,p222,p223);
FA fa69(ip_12_2,ip_13_1,ip_14_0,p224,p225);
HA ha43(p180,p184,p226,p227);
FA fa70(p215,p221,p223,p228,p229);
FA fa71(p190,p217,p219,p230,p231);
FA fa72(p225,p227,p182,p232,p233);
FA fa73(p186,p188,p194,p234,p235);
FA fa74(p229,p196,p198,p236,p237);
HA ha44(p231,p233,p238,p239);
FA fa75(p192,p235,p239,p240,p241);
HA ha45(p200,p237,p242,p243);
FA fa76(p202,p241,p243,p244,p245);
HA ha46(p204,p206,p246,p247);
HA ha47(p245,p247,p248,p249);
FA fa77(p208,p249,p210,p250,p251);
HA ha48(ip_0_15,ip_1_14,p252,p253);
HA ha49(ip_2_13,ip_3_12,p254,p255);
FA fa78(ip_4_11,ip_5_10,ip_6_9,p256,p257);
HA ha50(ip_7_8,ip_8_7,p258,p259);
HA ha51(ip_9_6,ip_10_5,p260,p261);
FA fa79(ip_11_4,ip_12_3,ip_13_2,p262,p263);
FA fa80(ip_14_1,ip_15_0,p214,p264,p265);
FA fa81(p220,p222,p253,p266,p267);
FA fa82(p255,p259,p261,p268,p269);
HA ha52(p226,p257,p270,p271);
FA fa83(p263,p265,p216,p272,p273);
FA fa84(p218,p224,p267,p274,p275);
FA fa85(p269,p271,p228,p276,p277);
FA fa86(p273,p230,p232,p278,p279);
HA ha53(p238,p275,p280,p281);
FA fa87(p277,p234,p281,p282,p283);
HA ha54(p236,p242,p284,p285);
FA fa88(p279,p240,p283,p286,p287);
HA ha55(p285,p244,p288,p289);
FA fa89(p246,p287,p248,p290,p291);
FA fa90(p289,p291,p250,p292,p293);
FA fa91(ip_1_15,ip_2_14,ip_3_13,p294,p295);
HA ha56(ip_4_12,ip_5_11,p296,p297);
HA ha57(ip_6_10,ip_7_9,p298,p299);
FA fa92(ip_8_8,ip_9_7,ip_10_6,p300,p301);
HA ha58(ip_11_5,ip_12_4,p302,p303);
FA fa93(ip_13_3,ip_14_2,ip_15_1,p304,p305);
HA ha59(p252,p254,p306,p307);
FA fa94(p258,p260,p297,p308,p309);
HA ha60(p299,p303,p310,p311);
HA ha61(p295,p301,p312,p313);
FA fa95(p305,p307,p311,p314,p315);
FA fa96(p256,p262,p264,p316,p317);
HA ha62(p270,p309,p318,p319);
HA ha63(p313,p266,p320,p321);
FA fa97(p268,p315,p319,p322,p323);
HA ha64(p272,p317,p324,p325);
HA ha65(p321,p274,p326,p327);
FA fa98(p276,p280,p323,p328,p329);
FA fa99(p325,p327,p278,p330,p331);
FA fa100(p284,p329,p282,p332,p333);
FA fa101(p331,p333,p286,p334,p335);
FA fa102(p288,p335,p290,p336,p337);
FA fa103(ip_2_15,ip_3_14,ip_4_13,p338,p339);
HA ha66(ip_5_12,ip_6_11,p340,p341);
FA fa104(ip_7_10,ip_8_9,ip_9_8,p342,p343);
HA ha67(ip_10_7,ip_11_6,p344,p345);
FA fa105(ip_12_5,ip_13_4,ip_14_3,p346,p347);
FA fa106(ip_15_2,p296,p298,p348,p349);
FA fa107(p302,p341,p345,p350,p351);
HA ha68(p306,p310,p352,p353);
FA fa108(p339,p343,p347,p354,p355);
FA fa109(p294,p300,p304,p356,p357);
FA fa110(p312,p349,p351,p358,p359);
FA fa111(p353,p308,p318,p360,p361);
HA ha69(p355,p314,p362,p363);
FA fa112(p320,p357,p359,p364,p365);
HA ha70(p316,p324,p366,p367);
HA ha71(p361,p363,p368,p369);
FA fa113(p322,p326,p365,p370,p371);
HA ha72(p367,p369,p372,p373);
HA ha73(p373,p328,p374,p375);
FA fa114(p371,p330,p375,p376,p377);
HA ha74(p332,p377,p378,p379);
HA ha75(p334,p379,p380,p381);
HA ha76(ip_3_15,ip_4_14,p382,p383);
HA ha77(ip_5_13,ip_6_12,p384,p385);
HA ha78(ip_7_11,ip_8_10,p386,p387);
FA fa115(ip_9_9,ip_10_8,ip_11_7,p388,p389);
FA fa116(ip_12_6,ip_13_5,ip_14_4,p390,p391);
HA ha79(ip_15_3,p340,p392,p393);
HA ha80(p344,p383,p394,p395);
HA ha81(p385,p387,p396,p397);
FA fa117(p389,p391,p393,p398,p399);
FA fa118(p395,p397,p338,p400,p401);
FA fa119(p342,p346,p352,p402,p403);
HA ha82(p348,p350,p404,p405);
HA ha83(p399,p401,p406,p407);
FA fa120(p354,p403,p405,p408,p409);
HA ha84(p407,p356,p410,p411);
FA fa121(p358,p362,p360,p412,p413);
HA ha85(p366,p368,p414,p415);
HA ha86(p409,p411,p416,p417);
FA fa122(p364,p372,p413,p418,p419);
FA fa123(p415,p417,p370,p420,p421);
FA fa124(p374,p419,p421,p422,p423);
HA ha87(p423,p376,p424,p425);
FA fa125(p378,p380,p425,p426,p427);
FA fa126(ip_4_15,ip_5_14,ip_6_13,p428,p429);
FA fa127(ip_7_12,ip_8_11,ip_9_10,p430,p431);
HA ha88(ip_10_9,ip_11_8,p432,p433);
FA fa128(ip_12_7,ip_13_6,ip_14_5,p434,p435);
FA fa129(ip_15_4,p382,p384,p436,p437);
FA fa130(p386,p433,p392,p438,p439);
FA fa131(p394,p396,p429,p440,p441);
FA fa132(p431,p435,p388,p442,p443);
FA fa133(p390,p437,p439,p444,p445);
FA fa134(p441,p443,p398,p446,p447);
HA ha89(p400,p404,p448,p449);
HA ha90(p406,p445,p450,p451);
HA ha91(p402,p447,p452,p453);
FA fa135(p449,p451,p410,p454,p455);
FA fa136(p453,p408,p414,p456,p457);
FA fa137(p416,p455,p412,p458,p459);
FA fa138(p457,p459,p418,p460,p461);
FA fa139(p420,p461,p422,p462,p463);
HA ha92(p424,p463,p464,p465);
HA ha93(ip_5_15,ip_6_14,p466,p467);
FA fa140(ip_7_13,ip_8_12,ip_9_11,p468,p469);
FA fa141(ip_10_10,ip_11_9,ip_12_8,p470,p471);
FA fa142(ip_13_7,ip_14_6,ip_15_5,p472,p473);
HA ha94(p432,p467,p474,p475);
FA fa143(p469,p471,p473,p476,p477);
FA fa144(p475,p428,p430,p478,p479);
FA fa145(p434,p436,p438,p480,p481);
HA ha95(p477,p440,p482,p483);
HA ha96(p442,p479,p484,p485);
FA fa146(p444,p448,p450,p486,p487);
HA ha97(p481,p483,p488,p489);
FA fa147(p485,p446,p452,p490,p491);
HA ha98(p489,p487,p492,p493);
FA fa148(p454,p491,p493,p494,p495);
FA fa149(p456,p458,p495,p496,p497);
FA fa150(p460,p497,p462,p498,p499);
HA ha99(ip_6_15,ip_7_14,p500,p501);
HA ha100(ip_8_13,ip_9_12,p502,p503);
HA ha101(ip_10_11,ip_11_10,p504,p505);
HA ha102(ip_12_9,ip_13_8,p506,p507);
HA ha103(ip_14_7,ip_15_6,p508,p509);
HA ha104(p466,p501,p510,p511);
FA fa151(p503,p505,p507,p512,p513);
FA fa152(p509,p474,p511,p514,p515);
HA ha105(p468,p470,p516,p517);
FA fa153(p472,p513,p515,p518,p519);
FA fa154(p517,p476,p519,p520,p521);
FA fa155(p478,p482,p484,p522,p523);
HA ha106(p480,p488,p524,p525);
FA fa156(p521,p523,p525,p526,p527);
FA fa157(p486,p492,p490,p528,p529);
HA ha107(p527,p529,p530,p531);
HA ha108(p494,p531,p532,p533);
FA fa158(p533,p496,p498,p534,p535);
HA ha109(ip_7_15,ip_8_14,p536,p537);
FA fa159(ip_9_13,ip_10_12,ip_11_11,p538,p539);
FA fa160(ip_12_10,ip_13_9,ip_14_8,p540,p541);
HA ha110(ip_15_7,p500,p542,p543);
HA ha111(p502,p504,p544,p545);
FA fa161(p506,p508,p537,p546,p547);
HA ha112(p510,p539,p548,p549);
HA ha113(p541,p543,p550,p551);
FA fa162(p545,p547,p549,p552,p553);
FA fa163(p551,p512,p516,p554,p555);
FA fa164(p514,p553,p518,p556,p557);
FA fa165(p555,p557,p520,p558,p559);
HA ha114(p524,p522,p560,p561);
HA ha115(p559,p561,p562,p563);
HA ha116(p526,p563,p564,p565);
HA ha117(p528,p530,p566,p567);
HA ha118(p565,p532,p568,p569);
HA ha119(p567,p569,p570,p571);
HA ha120(ip_8_15,ip_9_14,p572,p573);
HA ha121(ip_10_13,ip_11_12,p574,p575);
FA fa166(ip_12_11,ip_13_10,ip_14_9,p576,p577);
FA fa167(ip_15_8,p536,p573,p578,p579);
FA fa168(p575,p542,p544,p580,p581);
FA fa169(p577,p538,p540,p582,p583);
HA ha122(p548,p550,p584,p585);
HA ha123(p579,p546,p586,p587);
HA ha124(p581,p585,p588,p589);
FA fa170(p583,p587,p589,p590,p591);
HA ha125(p552,p554,p592,p593);
FA fa171(p591,p556,p593,p594,p595);
HA ha126(p558,p560,p596,p597);
HA ha127(p595,p562,p598,p599);
HA ha128(p597,p564,p600,p601);
FA fa172(p599,p566,p601,p602,p603);
HA ha129(p568,p570,p604,p605);
FA fa173(ip_9_15,ip_10_14,ip_11_13,p606,p607);
FA fa174(ip_12_12,ip_13_11,ip_14_10,p608,p609);
HA ha130(ip_15_9,p572,p610,p611);
FA fa175(p574,p607,p609,p612,p613);
HA ha131(p611,p576,p614,p615);
FA fa176(p578,p584,p613,p616,p617);
FA fa177(p615,p580,p586,p618,p619);
HA ha132(p588,p582,p620,p621);
FA fa178(p617,p619,p621,p622,p623);
HA ha133(p590,p592,p624,p625);
FA fa179(p623,p625,p594,p626,p627);
FA fa180(p596,p598,p627,p628,p629);
FA fa181(p600,p629,p602,p630,p631);
HA ha134(ip_10_15,ip_11_14,p632,p633);
HA ha135(ip_12_13,ip_13_12,p634,p635);
HA ha136(ip_14_11,ip_15_10,p636,p637);
HA ha137(p633,p635,p638,p639);
FA fa182(p637,p610,p639,p640,p641);
FA fa183(p606,p608,p614,p642,p643);
FA fa184(p641,p612,p643,p644,p645);
FA fa185(p616,p620,p645,p646,p647);
HA ha138(p618,p624,p648,p649);
FA fa186(p647,p622,p649,p650,p651);
HA ha139(p651,p626,p652,p653);
HA ha140(p653,p628,p654,p655);
HA ha141(ip_11_15,ip_12_14,p656,p657);
HA ha142(ip_13_13,ip_14_12,p658,p659);
FA fa187(ip_15_11,p632,p634,p660,p661);
HA ha143(p636,p657,p662,p663);
FA fa188(p659,p638,p663,p664,p665);
FA fa189(p661,p665,p640,p666,p667);
HA ha144(p642,p667,p668,p669);
FA fa190(p669,p644,p646,p670,p671);
HA ha145(p648,p671,p672,p673);
FA fa191(p673,p650,p652,p674,p675);
HA ha146(ip_12_15,ip_13_14,p676,p677);
HA ha147(ip_14_13,ip_15_12,p678,p679);
HA ha148(p656,p658,p680,p681);
HA ha149(p677,p679,p682,p683);
HA ha150(p662,p681,p684,p685);
FA fa192(p683,p685,p660,p686,p687);
FA fa193(p664,p687,p666,p688,p689);
FA fa194(p668,p689,p670,p690,p691);
HA ha151(p672,p691,p692,p693);
FA fa195(ip_13_15,ip_14_14,ip_15_13,p694,p695);
FA fa196(p676,p678,p680,p696,p697);
FA fa197(p682,p695,p684,p698,p699);
HA ha152(p697,p699,p700,p701);
FA fa198(p701,p686,p688,p702,p703);
HA ha153(p703,p690,p704,p705);
HA ha154(ip_14_15,ip_15_14,p706,p707);
HA ha155(p707,p694,p708,p709);
FA fa199(p696,p709,p698,p710,p711);
FA fa200(p700,p711,p702,p712,p713);
FA fa201(ip_15_15,p706,p708,p714,p715);
HA ha156(p715,p710,p716,p717);
wire [31:0] a,b;
wire [31:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p0;
assign b[3] = p5;
assign a[4] = p13;
assign b[4] = 1'b0;
assign a[5] = p12;
assign b[5] = p25;
assign a[6] = p24;
assign b[6] = p37;
assign a[7] = p53;
assign b[7] = 1'b0;
assign a[8] = p71;
assign b[8] = p52;
assign a[9] = p93;
assign b[9] = 1'b0;
assign a[10] = p117;
assign b[10] = 1'b0;
assign a[11] = p149;
assign b[11] = 1'b0;
assign a[12] = p179;
assign b[12] = p148;
assign a[13] = p213;
assign b[13] = p178;
assign a[14] = p212;
assign b[14] = p251;
assign a[15] = p293;
assign b[15] = 1'b0;
assign a[16] = p337;
assign b[16] = p292;
assign a[17] = p381;
assign b[17] = p336;
assign a[18] = p427;
assign b[18] = 1'b0;
assign a[19] = p465;
assign b[19] = p426;
assign a[20] = p464;
assign b[20] = p499;
assign a[21] = p535;
assign b[21] = 1'b0;
assign a[22] = p571;
assign b[22] = p534;
assign a[23] = p603;
assign b[23] = p605;
assign a[24] = p604;
assign b[24] = p631;
assign a[25] = p655;
assign b[25] = p630;
assign a[26] = p675;
assign b[26] = p654;
assign a[27] = p693;
assign b[27] = p674;
assign a[28] = p692;
assign b[28] = p705;
assign a[29] = p713;
assign b[29] = p704;
assign a[30] = p717;
assign b[30] = p712;
assign a[31] = p714;
assign b[31] = p716;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[31] = s[31];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [31:0] a,b;
output [31:0] s;
assign s = a+b;
endmodule
