// 1 2 2 2 2 2 2 2 2 1 1 2 1 2 1 2 

module main(x,y,o);
input [7:0] x,y;
output [15:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_1_0,x[1],y[0]);
and and9(ip_1_1,x[1],y[1]);
and and10(ip_1_2,x[1],y[2]);
and and11(ip_1_3,x[1],y[3]);
and and12(ip_1_4,x[1],y[4]);
and and13(ip_1_5,x[1],y[5]);
and and14(ip_1_6,x[1],y[6]);
and and15(ip_1_7,x[1],y[7]);
and and16(ip_2_0,x[2],y[0]);
and and17(ip_2_1,x[2],y[1]);
and and18(ip_2_2,x[2],y[2]);
and and19(ip_2_3,x[2],y[3]);
and and20(ip_2_4,x[2],y[4]);
and and21(ip_2_5,x[2],y[5]);
and and22(ip_2_6,x[2],y[6]);
and and23(ip_2_7,x[2],y[7]);
and and24(ip_3_0,x[3],y[0]);
and and25(ip_3_1,x[3],y[1]);
and and26(ip_3_2,x[3],y[2]);
and and27(ip_3_3,x[3],y[3]);
and and28(ip_3_4,x[3],y[4]);
and and29(ip_3_5,x[3],y[5]);
and and30(ip_3_6,x[3],y[6]);
and and31(ip_3_7,x[3],y[7]);
and and32(ip_4_0,x[4],y[0]);
and and33(ip_4_1,x[4],y[1]);
and and34(ip_4_2,x[4],y[2]);
and and35(ip_4_3,x[4],y[3]);
and and36(ip_4_4,x[4],y[4]);
and and37(ip_4_5,x[4],y[5]);
and and38(ip_4_6,x[4],y[6]);
and and39(ip_4_7,x[4],y[7]);
and and40(ip_5_0,x[5],y[0]);
and and41(ip_5_1,x[5],y[1]);
and and42(ip_5_2,x[5],y[2]);
and and43(ip_5_3,x[5],y[3]);
and and44(ip_5_4,x[5],y[4]);
and and45(ip_5_5,x[5],y[5]);
and and46(ip_5_6,x[5],y[6]);
and and47(ip_5_7,x[5],y[7]);
and and48(ip_6_0,x[6],y[0]);
and and49(ip_6_1,x[6],y[1]);
and and50(ip_6_2,x[6],y[2]);
and and51(ip_6_3,x[6],y[3]);
and and52(ip_6_4,x[6],y[4]);
and and53(ip_6_5,x[6],y[5]);
and and54(ip_6_6,x[6],y[6]);
and and55(ip_6_7,x[6],y[7]);
and and56(ip_7_0,x[7],y[0]);
and and57(ip_7_1,x[7],y[1]);
and and58(ip_7_2,x[7],y[2]);
and and59(ip_7_3,x[7],y[3]);
and and60(ip_7_4,x[7],y[4]);
and and61(ip_7_5,x[7],y[5]);
and and62(ip_7_6,x[7],y[6]);
and and63(ip_7_7,x[7],y[7]);
HA ha0(ip_0_2,ip_1_1,p0,p1);
HA ha1(ip_0_3,ip_1_2,p2,p3);
FA fa0(ip_2_1,ip_3_0,p0,p4,p5);
HA ha2(ip_0_4,ip_1_3,p6,p7);
HA ha3(ip_2_2,ip_3_1,p8,p9);
HA ha4(ip_4_0,p2,p10,p11);
HA ha5(p7,p9,p12,p13);
HA ha6(p11,p13,p14,p15);
FA fa1(ip_0_5,ip_1_4,ip_2_3,p16,p17);
HA ha7(ip_3_2,ip_4_1,p18,p19);
FA fa2(ip_5_0,p19,p6,p20,p21);
HA ha8(p8,p10,p22,p23);
FA fa3(p12,p17,p14,p24,p25);
HA ha9(p21,p23,p26,p27);
HA ha10(ip_0_6,ip_1_5,p28,p29);
FA fa4(ip_2_4,ip_3_3,ip_4_2,p30,p31);
FA fa5(ip_5_1,ip_6_0,p18,p32,p33);
HA ha11(p29,p31,p34,p35);
HA ha12(p33,p16,p36,p37);
FA fa6(p22,p35,p20,p38,p39);
FA fa7(p26,p37,p24,p40,p41);
HA ha13(ip_0_7,ip_1_6,p42,p43);
HA ha14(ip_2_5,ip_3_4,p44,p45);
FA fa8(ip_4_3,ip_5_2,ip_6_1,p46,p47);
FA fa9(ip_7_0,p28,p43,p48,p49);
FA fa10(p45,p47,p30,p50,p51);
FA fa11(p32,p34,p49,p52,p53);
FA fa12(p36,p51,p53,p54,p55);
HA ha15(p38,p55,p56,p57);
HA ha16(ip_1_7,ip_2_6,p58,p59);
FA fa13(ip_3_5,ip_4_4,ip_5_3,p60,p61);
HA ha17(ip_6_2,ip_7_1,p62,p63);
HA ha18(p42,p44,p64,p65);
FA fa14(p59,p63,p61,p66,p67);
HA ha19(p65,p46,p68,p69);
HA ha20(p67,p48,p70,p71);
HA ha21(p69,p50,p72,p73);
HA ha22(p71,p52,p74,p75);
HA ha23(p73,p54,p76,p77);
HA ha24(p56,p75,p78,p79);
HA ha25(ip_2_7,ip_3_6,p80,p81);
FA fa15(ip_4_5,ip_5_4,ip_6_3,p82,p83);
HA ha26(ip_7_2,p58,p84,p85);
FA fa16(p62,p81,p64,p86,p87);
FA fa17(p83,p85,p60,p88,p89);
FA fa18(p87,p66,p68,p90,p91);
FA fa19(p89,p70,p72,p92,p93);
HA ha27(p91,p74,p94,p95);
HA ha28(p93,p76,p96,p97);
FA fa20(p78,p95,p97,p98,p99);
HA ha29(ip_3_7,ip_4_6,p100,p101);
FA fa21(ip_5_5,ip_6_4,ip_7_3,p102,p103);
HA ha30(p101,p80,p104,p105);
FA fa22(p103,p105,p84,p106,p107);
FA fa23(p82,p107,p86,p108,p109);
FA fa24(p88,p109,p90,p110,p111);
FA fa25(p111,p92,p94,p112,p113);
FA fa26(p96,p113,p98,p114,p115);
FA fa27(ip_4_7,ip_5_6,ip_6_5,p116,p117);
FA fa28(ip_7_4,p100,p104,p118,p119);
FA fa29(p117,p102,p119,p120,p121);
HA ha31(p106,p121,p122,p123);
FA fa30(p123,p108,p110,p124,p125);
HA ha32(p125,p112,p126,p127);
FA fa31(ip_5_7,ip_6_6,ip_7_5,p128,p129);
FA fa32(p129,p116,p118,p130,p131);
HA ha33(p131,p120,p132,p133);
HA ha34(p122,p133,p134,p135);
FA fa33(p135,p124,p126,p136,p137);
FA fa34(ip_6_7,ip_7_6,p128,p138,p139);
HA ha35(p139,p130,p140,p141);
FA fa35(p132,p141,p134,p142,p143);
HA ha36(ip_7_7,p138,p144,p145);
FA fa36(p145,p140,p142,p146,p147);
wire [15:0] a,b;
wire [15:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = ip_2_0;
assign b[2] = p1;
assign a[3] = p3;
assign b[3] = p5;
assign a[4] = p15;
assign b[4] = p4;
assign a[5] = p25;
assign b[5] = p27;
assign a[6] = p39;
assign b[6] = p41;
assign a[7] = p40;
assign b[7] = p57;
assign a[8] = p77;
assign b[8] = p79;
assign a[9] = p99;
assign b[9] = 1'b0;
assign a[10] = p115;
assign b[10] = 1'b0;
assign a[11] = p127;
assign b[11] = p114;
assign a[12] = p137;
assign b[12] = 1'b0;
assign a[13] = p143;
assign b[13] = p136;
assign a[14] = p147;
assign b[14] = 1'b0;
assign a[15] = p144;
assign b[15] = p146;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[15] = s[15];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [15:0] a,b;
output [15:0] s;
assign s = a+b;
endmodule
