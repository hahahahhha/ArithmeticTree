// 1 2 1 1 1 2 1 2 1 2 2 2 2 2 2 1 1 1 1 1 2 1 2 2 

module main(x,y,o);
input [11:0] x,y;
output [23:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_1_0,x[1],y[0]);
and and13(ip_1_1,x[1],y[1]);
and and14(ip_1_2,x[1],y[2]);
and and15(ip_1_3,x[1],y[3]);
and and16(ip_1_4,x[1],y[4]);
and and17(ip_1_5,x[1],y[5]);
and and18(ip_1_6,x[1],y[6]);
and and19(ip_1_7,x[1],y[7]);
and and20(ip_1_8,x[1],y[8]);
and and21(ip_1_9,x[1],y[9]);
and and22(ip_1_10,x[1],y[10]);
and and23(ip_1_11,x[1],y[11]);
and and24(ip_2_0,x[2],y[0]);
and and25(ip_2_1,x[2],y[1]);
and and26(ip_2_2,x[2],y[2]);
and and27(ip_2_3,x[2],y[3]);
and and28(ip_2_4,x[2],y[4]);
and and29(ip_2_5,x[2],y[5]);
and and30(ip_2_6,x[2],y[6]);
and and31(ip_2_7,x[2],y[7]);
and and32(ip_2_8,x[2],y[8]);
and and33(ip_2_9,x[2],y[9]);
and and34(ip_2_10,x[2],y[10]);
and and35(ip_2_11,x[2],y[11]);
and and36(ip_3_0,x[3],y[0]);
and and37(ip_3_1,x[3],y[1]);
and and38(ip_3_2,x[3],y[2]);
and and39(ip_3_3,x[3],y[3]);
and and40(ip_3_4,x[3],y[4]);
and and41(ip_3_5,x[3],y[5]);
and and42(ip_3_6,x[3],y[6]);
and and43(ip_3_7,x[3],y[7]);
and and44(ip_3_8,x[3],y[8]);
and and45(ip_3_9,x[3],y[9]);
and and46(ip_3_10,x[3],y[10]);
and and47(ip_3_11,x[3],y[11]);
and and48(ip_4_0,x[4],y[0]);
and and49(ip_4_1,x[4],y[1]);
and and50(ip_4_2,x[4],y[2]);
and and51(ip_4_3,x[4],y[3]);
and and52(ip_4_4,x[4],y[4]);
and and53(ip_4_5,x[4],y[5]);
and and54(ip_4_6,x[4],y[6]);
and and55(ip_4_7,x[4],y[7]);
and and56(ip_4_8,x[4],y[8]);
and and57(ip_4_9,x[4],y[9]);
and and58(ip_4_10,x[4],y[10]);
and and59(ip_4_11,x[4],y[11]);
and and60(ip_5_0,x[5],y[0]);
and and61(ip_5_1,x[5],y[1]);
and and62(ip_5_2,x[5],y[2]);
and and63(ip_5_3,x[5],y[3]);
and and64(ip_5_4,x[5],y[4]);
and and65(ip_5_5,x[5],y[5]);
and and66(ip_5_6,x[5],y[6]);
and and67(ip_5_7,x[5],y[7]);
and and68(ip_5_8,x[5],y[8]);
and and69(ip_5_9,x[5],y[9]);
and and70(ip_5_10,x[5],y[10]);
and and71(ip_5_11,x[5],y[11]);
and and72(ip_6_0,x[6],y[0]);
and and73(ip_6_1,x[6],y[1]);
and and74(ip_6_2,x[6],y[2]);
and and75(ip_6_3,x[6],y[3]);
and and76(ip_6_4,x[6],y[4]);
and and77(ip_6_5,x[6],y[5]);
and and78(ip_6_6,x[6],y[6]);
and and79(ip_6_7,x[6],y[7]);
and and80(ip_6_8,x[6],y[8]);
and and81(ip_6_9,x[6],y[9]);
and and82(ip_6_10,x[6],y[10]);
and and83(ip_6_11,x[6],y[11]);
and and84(ip_7_0,x[7],y[0]);
and and85(ip_7_1,x[7],y[1]);
and and86(ip_7_2,x[7],y[2]);
and and87(ip_7_3,x[7],y[3]);
and and88(ip_7_4,x[7],y[4]);
and and89(ip_7_5,x[7],y[5]);
and and90(ip_7_6,x[7],y[6]);
and and91(ip_7_7,x[7],y[7]);
and and92(ip_7_8,x[7],y[8]);
and and93(ip_7_9,x[7],y[9]);
and and94(ip_7_10,x[7],y[10]);
and and95(ip_7_11,x[7],y[11]);
and and96(ip_8_0,x[8],y[0]);
and and97(ip_8_1,x[8],y[1]);
and and98(ip_8_2,x[8],y[2]);
and and99(ip_8_3,x[8],y[3]);
and and100(ip_8_4,x[8],y[4]);
and and101(ip_8_5,x[8],y[5]);
and and102(ip_8_6,x[8],y[6]);
and and103(ip_8_7,x[8],y[7]);
and and104(ip_8_8,x[8],y[8]);
and and105(ip_8_9,x[8],y[9]);
and and106(ip_8_10,x[8],y[10]);
and and107(ip_8_11,x[8],y[11]);
and and108(ip_9_0,x[9],y[0]);
and and109(ip_9_1,x[9],y[1]);
and and110(ip_9_2,x[9],y[2]);
and and111(ip_9_3,x[9],y[3]);
and and112(ip_9_4,x[9],y[4]);
and and113(ip_9_5,x[9],y[5]);
and and114(ip_9_6,x[9],y[6]);
and and115(ip_9_7,x[9],y[7]);
and and116(ip_9_8,x[9],y[8]);
and and117(ip_9_9,x[9],y[9]);
and and118(ip_9_10,x[9],y[10]);
and and119(ip_9_11,x[9],y[11]);
and and120(ip_10_0,x[10],y[0]);
and and121(ip_10_1,x[10],y[1]);
and and122(ip_10_2,x[10],y[2]);
and and123(ip_10_3,x[10],y[3]);
and and124(ip_10_4,x[10],y[4]);
and and125(ip_10_5,x[10],y[5]);
and and126(ip_10_6,x[10],y[6]);
and and127(ip_10_7,x[10],y[7]);
and and128(ip_10_8,x[10],y[8]);
and and129(ip_10_9,x[10],y[9]);
and and130(ip_10_10,x[10],y[10]);
and and131(ip_10_11,x[10],y[11]);
and and132(ip_11_0,x[11],y[0]);
and and133(ip_11_1,x[11],y[1]);
and and134(ip_11_2,x[11],y[2]);
and and135(ip_11_3,x[11],y[3]);
and and136(ip_11_4,x[11],y[4]);
and and137(ip_11_5,x[11],y[5]);
and and138(ip_11_6,x[11],y[6]);
and and139(ip_11_7,x[11],y[7]);
and and140(ip_11_8,x[11],y[8]);
and and141(ip_11_9,x[11],y[9]);
and and142(ip_11_10,x[11],y[10]);
and and143(ip_11_11,x[11],y[11]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
FA fa2(ip_3_0,p3,p0,p4,p5);
HA ha0(ip_0_4,ip_1_3,p6,p7);
FA fa3(ip_2_2,ip_3_1,ip_4_0,p8,p9);
HA ha1(p7,p9,p10,p11);
FA fa4(p11,p2,p4,p12,p13);
HA ha2(ip_0_5,ip_1_4,p14,p15);
HA ha3(ip_2_3,ip_3_2,p16,p17);
FA fa5(ip_4_1,ip_5_0,p15,p18,p19);
HA ha4(p17,p6,p20,p21);
HA ha5(p19,p21,p22,p23);
HA ha6(p10,p23,p24,p25);
HA ha7(p8,p25,p26,p27);
FA fa6(ip_0_6,ip_1_5,ip_2_4,p28,p29);
FA fa7(ip_3_3,ip_4_2,ip_5_1,p30,p31);
FA fa8(ip_6_0,p14,p16,p32,p33);
HA ha8(p20,p29,p34,p35);
FA fa9(p31,p18,p22,p36,p37);
FA fa10(p33,p35,p24,p38,p39);
FA fa11(p26,p37,p39,p40,p41);
FA fa12(ip_0_7,ip_1_6,ip_2_5,p42,p43);
FA fa13(ip_3_4,ip_4_3,ip_5_2,p44,p45);
FA fa14(ip_6_1,ip_7_0,p43,p46,p47);
FA fa15(p45,p28,p30,p48,p49);
FA fa16(p34,p47,p32,p50,p51);
HA ha9(p49,p51,p52,p53);
FA fa17(p36,p38,p53,p54,p55);
HA ha10(ip_0_8,ip_1_7,p56,p57);
FA fa18(ip_2_6,ip_3_5,ip_4_4,p58,p59);
HA ha11(ip_5_3,ip_6_2,p60,p61);
HA ha12(ip_7_1,ip_8_0,p62,p63);
FA fa19(p57,p61,p63,p64,p65);
FA fa20(p59,p42,p44,p66,p67);
FA fa21(p65,p46,p67,p68,p69);
FA fa22(p48,p50,p52,p70,p71);
FA fa23(p69,p71,p54,p72,p73);
FA fa24(ip_0_9,ip_1_8,ip_2_7,p74,p75);
FA fa25(ip_3_6,ip_4_5,ip_5_4,p76,p77);
FA fa26(ip_6_3,ip_7_2,ip_8_1,p78,p79);
FA fa27(ip_9_0,p56,p60,p80,p81);
HA ha13(p62,p75,p82,p83);
HA ha14(p77,p79,p84,p85);
FA fa28(p58,p81,p83,p86,p87);
HA ha15(p85,p64,p88,p89);
HA ha16(p87,p89,p90,p91);
HA ha17(p66,p91,p92,p93);
FA fa29(p68,p93,p70,p94,p95);
FA fa30(ip_0_10,ip_1_9,ip_2_8,p96,p97);
FA fa31(ip_3_7,ip_4_6,ip_5_5,p98,p99);
HA ha18(ip_6_4,ip_7_3,p100,p101);
FA fa32(ip_8_2,ip_9_1,ip_10_0,p102,p103);
HA ha19(p101,p103,p104,p105);
HA ha20(p97,p99,p106,p107);
FA fa33(p105,p107,p74,p108,p109);
HA ha21(p76,p78,p110,p111);
FA fa34(p82,p84,p111,p112,p113);
HA ha22(p80,p109,p114,p115);
HA ha23(p113,p88,p116,p117);
HA ha24(p115,p117,p118,p119);
HA ha25(p86,p90,p120,p121);
FA fa35(p119,p121,p92,p122,p123);
FA fa36(ip_0_11,ip_1_10,ip_2_9,p124,p125);
FA fa37(ip_3_8,ip_4_7,ip_5_6,p126,p127);
HA ha26(ip_6_5,ip_7_4,p128,p129);
HA ha27(ip_8_3,ip_9_2,p130,p131);
HA ha28(ip_10_1,ip_11_0,p132,p133);
FA fa38(p100,p129,p131,p134,p135);
FA fa39(p133,p125,p127,p136,p137);
HA ha29(p102,p104,p138,p139);
FA fa40(p106,p135,p96,p140,p141);
HA ha30(p98,p110,p142,p143);
FA fa41(p137,p139,p141,p144,p145);
HA ha31(p143,p108,p146,p147);
FA fa42(p112,p114,p116,p148,p149);
FA fa43(p145,p118,p120,p150,p151);
FA fa44(p147,p149,p151,p152,p153);
FA fa45(ip_1_11,ip_2_10,ip_3_9,p154,p155);
HA ha32(ip_4_8,ip_5_7,p156,p157);
HA ha33(ip_6_6,ip_7_5,p158,p159);
HA ha34(ip_8_4,ip_9_3,p160,p161);
FA fa46(ip_10_2,ip_11_1,p128,p162,p163);
FA fa47(p130,p132,p157,p164,p165);
FA fa48(p159,p161,p155,p166,p167);
HA ha35(p163,p124,p168,p169);
FA fa49(p126,p165,p167,p170,p171);
HA ha36(p134,p138,p172,p173);
FA fa50(p169,p136,p142,p174,p175);
FA fa51(p171,p173,p140,p176,p177);
HA ha37(p144,p146,p178,p179);
FA fa52(p175,p177,p179,p180,p181);
HA ha38(p148,p181,p182,p183);
HA ha39(p150,p183,p184,p185);
HA ha40(ip_2_11,ip_3_10,p186,p187);
HA ha41(ip_4_9,ip_5_8,p188,p189);
HA ha42(ip_6_7,ip_7_6,p190,p191);
FA fa53(ip_8_5,ip_9_4,ip_10_3,p192,p193);
FA fa54(ip_11_2,p156,p158,p194,p195);
HA ha43(p160,p187,p196,p197);
FA fa55(p189,p191,p193,p198,p199);
FA fa56(p197,p154,p162,p200,p201);
HA ha44(p195,p199,p202,p203);
FA fa57(p164,p166,p168,p204,p205);
HA ha45(p203,p172,p206,p207);
HA ha46(p201,p170,p208,p209);
HA ha47(p205,p207,p210,p211);
FA fa58(p209,p211,p174,p212,p213);
FA fa59(p176,p178,p213,p214,p215);
FA fa60(p180,p182,p215,p216,p217);
FA fa61(ip_3_11,ip_4_10,ip_5_9,p218,p219);
FA fa62(ip_6_8,ip_7_7,ip_8_6,p220,p221);
FA fa63(ip_9_5,ip_10_4,ip_11_3,p222,p223);
FA fa64(p186,p188,p190,p224,p225);
HA ha48(p196,p219,p226,p227);
HA ha49(p221,p223,p228,p229);
HA ha50(p192,p225,p230,p231);
FA fa65(p227,p229,p194,p232,p233);
FA fa66(p198,p202,p231,p234,p235);
HA ha51(p233,p200,p236,p237);
FA fa67(p206,p235,p204,p238,p239);
HA ha52(p208,p210,p240,p241);
FA fa68(p237,p239,p241,p242,p243);
FA fa69(p212,p243,p214,p244,p245);
FA fa70(ip_4_11,ip_5_10,ip_6_9,p246,p247);
HA ha53(ip_7_8,ip_8_7,p248,p249);
FA fa71(ip_9_6,ip_10_5,ip_11_4,p250,p251);
FA fa72(p249,p247,p251,p252,p253);
HA ha54(p218,p220,p254,p255);
FA fa73(p222,p226,p228,p256,p257);
FA fa74(p224,p230,p253,p258,p259);
FA fa75(p255,p257,p232,p260,p261);
FA fa76(p259,p234,p236,p262,p263);
FA fa77(p261,p240,p238,p264,p265);
HA ha55(p263,p265,p266,p267);
FA fa78(p242,p267,p244,p268,p269);
FA fa79(ip_5_11,ip_6_10,ip_7_9,p270,p271);
HA ha56(ip_8_8,ip_9_7,p272,p273);
HA ha57(ip_10_6,ip_11_5,p274,p275);
HA ha58(p248,p273,p276,p277);
FA fa80(p275,p271,p277,p278,p279);
HA ha59(p246,p250,p280,p281);
HA ha60(p254,p279,p282,p283);
HA ha61(p281,p252,p284,p285);
FA fa81(p283,p256,p285,p286,p287);
FA fa82(p258,p260,p287,p288,p289);
FA fa83(p262,p289,p264,p290,p291);
FA fa84(p266,p291,p268,p292,p293);
FA fa85(ip_6_11,ip_7_10,ip_8_9,p294,p295);
HA ha62(ip_9_8,ip_10_7,p296,p297);
FA fa86(ip_11_6,p272,p274,p298,p299);
HA ha63(p297,p276,p300,p301);
HA ha64(p295,p270,p302,p303);
FA fa87(p299,p301,p280,p304,p305);
HA ha65(p303,p278,p306,p307);
HA ha66(p282,p305,p308,p309);
FA fa88(p284,p307,p309,p310,p311);
HA ha67(p311,p286,p312,p313);
HA ha68(p313,p288,p314,p315);
FA fa89(p315,p290,p292,p316,p317);
HA ha69(ip_7_11,ip_8_10,p318,p319);
HA ha70(ip_9_9,ip_10_8,p320,p321);
FA fa90(ip_11_7,p296,p319,p322,p323);
FA fa91(p321,p294,p300,p324,p325);
FA fa92(p323,p298,p302,p326,p327);
FA fa93(p325,p304,p306,p328,p329);
FA fa94(p308,p327,p329,p330,p331);
FA fa95(p310,p331,p312,p332,p333);
FA fa96(p333,p314,p316,p334,p335);
FA fa97(ip_8_11,ip_9_10,ip_10_9,p336,p337);
HA ha71(ip_11_8,p318,p338,p339);
HA ha72(p320,p337,p340,p341);
HA ha73(p339,p341,p342,p343);
HA ha74(p322,p343,p344,p345);
HA ha75(p345,p324,p346,p347);
HA ha76(p326,p347,p348,p349);
FA fa98(p349,p328,p330,p350,p351);
FA fa99(p351,p332,p334,p352,p353);
FA fa100(ip_9_11,ip_10_10,ip_11_9,p354,p355);
HA ha77(p338,p355,p356,p357);
FA fa101(p336,p340,p357,p358,p359);
FA fa102(p342,p344,p359,p360,p361);
HA ha78(p346,p361,p362,p363);
FA fa103(p348,p363,p350,p364,p365);
FA fa104(ip_10_11,ip_11_10,p354,p366,p367);
FA fa105(p356,p367,p358,p368,p369);
HA ha79(p369,p360,p370,p371);
FA fa106(p362,p371,p364,p372,p373);
HA ha80(ip_11_11,p366,p374,p375);
FA fa107(p375,p368,p370,p376,p377);
wire [23:0] a,b;
wire [23:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p5;
assign b[3] = 1'b0;
assign a[4] = p13;
assign b[4] = 1'b0;
assign a[5] = p27;
assign b[5] = p12;
assign a[6] = p41;
assign b[6] = 1'b0;
assign a[7] = p40;
assign b[7] = p55;
assign a[8] = p73;
assign b[8] = 1'b0;
assign a[9] = p95;
assign b[9] = p72;
assign a[10] = p123;
assign b[10] = p94;
assign a[11] = p122;
assign b[11] = p153;
assign a[12] = p152;
assign b[12] = p185;
assign a[13] = p184;
assign b[13] = p217;
assign a[14] = p245;
assign b[14] = p216;
assign a[15] = p269;
assign b[15] = 1'b0;
assign a[16] = p293;
assign b[16] = 1'b0;
assign a[17] = p317;
assign b[17] = 1'b0;
assign a[18] = p335;
assign b[18] = 1'b0;
assign a[19] = p353;
assign b[19] = 1'b0;
assign a[20] = p365;
assign b[20] = p352;
assign a[21] = p373;
assign b[21] = 1'b0;
assign a[22] = p377;
assign b[22] = p372;
assign a[23] = p374;
assign b[23] = p376;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[23] = s[23];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [23:0] a,b;
output [23:0] s;
assign s = a+b;
endmodule
