// 1 2 1 2 2 1 2 2 2 1 2 2 2 2 2 2 1 1 1 2 2 2 1 2 2 1 2 2 2 2 2 1 2 2 1 2 2 2 2 2 2 2 2 1 2 2 1 2 1 1 2 2 2 2 2 2 2 1 2 2 2 1 2 3 

module main(x,y,o);
input [31:0] x,y;
output [63:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_0_16,ip_0_17,ip_0_18,ip_0_19,ip_0_20,ip_0_21,ip_0_22,ip_0_23,ip_0_24,ip_0_25,ip_0_26,ip_0_27,ip_0_28,ip_0_29,ip_0_30,ip_0_31,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_1_16,ip_1_17,ip_1_18,ip_1_19,ip_1_20,ip_1_21,ip_1_22,ip_1_23,ip_1_24,ip_1_25,ip_1_26,ip_1_27,ip_1_28,ip_1_29,ip_1_30,ip_1_31,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_2_16,ip_2_17,ip_2_18,ip_2_19,ip_2_20,ip_2_21,ip_2_22,ip_2_23,ip_2_24,ip_2_25,ip_2_26,ip_2_27,ip_2_28,ip_2_29,ip_2_30,ip_2_31,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_3_16,ip_3_17,ip_3_18,ip_3_19,ip_3_20,ip_3_21,ip_3_22,ip_3_23,ip_3_24,ip_3_25,ip_3_26,ip_3_27,ip_3_28,ip_3_29,ip_3_30,ip_3_31,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_4_16,ip_4_17,ip_4_18,ip_4_19,ip_4_20,ip_4_21,ip_4_22,ip_4_23,ip_4_24,ip_4_25,ip_4_26,ip_4_27,ip_4_28,ip_4_29,ip_4_30,ip_4_31,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_5_16,ip_5_17,ip_5_18,ip_5_19,ip_5_20,ip_5_21,ip_5_22,ip_5_23,ip_5_24,ip_5_25,ip_5_26,ip_5_27,ip_5_28,ip_5_29,ip_5_30,ip_5_31,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_6_16,ip_6_17,ip_6_18,ip_6_19,ip_6_20,ip_6_21,ip_6_22,ip_6_23,ip_6_24,ip_6_25,ip_6_26,ip_6_27,ip_6_28,ip_6_29,ip_6_30,ip_6_31,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_7_16,ip_7_17,ip_7_18,ip_7_19,ip_7_20,ip_7_21,ip_7_22,ip_7_23,ip_7_24,ip_7_25,ip_7_26,ip_7_27,ip_7_28,ip_7_29,ip_7_30,ip_7_31,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_8_16,ip_8_17,ip_8_18,ip_8_19,ip_8_20,ip_8_21,ip_8_22,ip_8_23,ip_8_24,ip_8_25,ip_8_26,ip_8_27,ip_8_28,ip_8_29,ip_8_30,ip_8_31,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_9_16,ip_9_17,ip_9_18,ip_9_19,ip_9_20,ip_9_21,ip_9_22,ip_9_23,ip_9_24,ip_9_25,ip_9_26,ip_9_27,ip_9_28,ip_9_29,ip_9_30,ip_9_31,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_10_16,ip_10_17,ip_10_18,ip_10_19,ip_10_20,ip_10_21,ip_10_22,ip_10_23,ip_10_24,ip_10_25,ip_10_26,ip_10_27,ip_10_28,ip_10_29,ip_10_30,ip_10_31,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_11_16,ip_11_17,ip_11_18,ip_11_19,ip_11_20,ip_11_21,ip_11_22,ip_11_23,ip_11_24,ip_11_25,ip_11_26,ip_11_27,ip_11_28,ip_11_29,ip_11_30,ip_11_31,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_12_16,ip_12_17,ip_12_18,ip_12_19,ip_12_20,ip_12_21,ip_12_22,ip_12_23,ip_12_24,ip_12_25,ip_12_26,ip_12_27,ip_12_28,ip_12_29,ip_12_30,ip_12_31,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_13_16,ip_13_17,ip_13_18,ip_13_19,ip_13_20,ip_13_21,ip_13_22,ip_13_23,ip_13_24,ip_13_25,ip_13_26,ip_13_27,ip_13_28,ip_13_29,ip_13_30,ip_13_31,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_14_16,ip_14_17,ip_14_18,ip_14_19,ip_14_20,ip_14_21,ip_14_22,ip_14_23,ip_14_24,ip_14_25,ip_14_26,ip_14_27,ip_14_28,ip_14_29,ip_14_30,ip_14_31,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15,ip_15_16,ip_15_17,ip_15_18,ip_15_19,ip_15_20,ip_15_21,ip_15_22,ip_15_23,ip_15_24,ip_15_25,ip_15_26,ip_15_27,ip_15_28,ip_15_29,ip_15_30,ip_15_31,ip_16_0,ip_16_1,ip_16_2,ip_16_3,ip_16_4,ip_16_5,ip_16_6,ip_16_7,ip_16_8,ip_16_9,ip_16_10,ip_16_11,ip_16_12,ip_16_13,ip_16_14,ip_16_15,ip_16_16,ip_16_17,ip_16_18,ip_16_19,ip_16_20,ip_16_21,ip_16_22,ip_16_23,ip_16_24,ip_16_25,ip_16_26,ip_16_27,ip_16_28,ip_16_29,ip_16_30,ip_16_31,ip_17_0,ip_17_1,ip_17_2,ip_17_3,ip_17_4,ip_17_5,ip_17_6,ip_17_7,ip_17_8,ip_17_9,ip_17_10,ip_17_11,ip_17_12,ip_17_13,ip_17_14,ip_17_15,ip_17_16,ip_17_17,ip_17_18,ip_17_19,ip_17_20,ip_17_21,ip_17_22,ip_17_23,ip_17_24,ip_17_25,ip_17_26,ip_17_27,ip_17_28,ip_17_29,ip_17_30,ip_17_31,ip_18_0,ip_18_1,ip_18_2,ip_18_3,ip_18_4,ip_18_5,ip_18_6,ip_18_7,ip_18_8,ip_18_9,ip_18_10,ip_18_11,ip_18_12,ip_18_13,ip_18_14,ip_18_15,ip_18_16,ip_18_17,ip_18_18,ip_18_19,ip_18_20,ip_18_21,ip_18_22,ip_18_23,ip_18_24,ip_18_25,ip_18_26,ip_18_27,ip_18_28,ip_18_29,ip_18_30,ip_18_31,ip_19_0,ip_19_1,ip_19_2,ip_19_3,ip_19_4,ip_19_5,ip_19_6,ip_19_7,ip_19_8,ip_19_9,ip_19_10,ip_19_11,ip_19_12,ip_19_13,ip_19_14,ip_19_15,ip_19_16,ip_19_17,ip_19_18,ip_19_19,ip_19_20,ip_19_21,ip_19_22,ip_19_23,ip_19_24,ip_19_25,ip_19_26,ip_19_27,ip_19_28,ip_19_29,ip_19_30,ip_19_31,ip_20_0,ip_20_1,ip_20_2,ip_20_3,ip_20_4,ip_20_5,ip_20_6,ip_20_7,ip_20_8,ip_20_9,ip_20_10,ip_20_11,ip_20_12,ip_20_13,ip_20_14,ip_20_15,ip_20_16,ip_20_17,ip_20_18,ip_20_19,ip_20_20,ip_20_21,ip_20_22,ip_20_23,ip_20_24,ip_20_25,ip_20_26,ip_20_27,ip_20_28,ip_20_29,ip_20_30,ip_20_31,ip_21_0,ip_21_1,ip_21_2,ip_21_3,ip_21_4,ip_21_5,ip_21_6,ip_21_7,ip_21_8,ip_21_9,ip_21_10,ip_21_11,ip_21_12,ip_21_13,ip_21_14,ip_21_15,ip_21_16,ip_21_17,ip_21_18,ip_21_19,ip_21_20,ip_21_21,ip_21_22,ip_21_23,ip_21_24,ip_21_25,ip_21_26,ip_21_27,ip_21_28,ip_21_29,ip_21_30,ip_21_31,ip_22_0,ip_22_1,ip_22_2,ip_22_3,ip_22_4,ip_22_5,ip_22_6,ip_22_7,ip_22_8,ip_22_9,ip_22_10,ip_22_11,ip_22_12,ip_22_13,ip_22_14,ip_22_15,ip_22_16,ip_22_17,ip_22_18,ip_22_19,ip_22_20,ip_22_21,ip_22_22,ip_22_23,ip_22_24,ip_22_25,ip_22_26,ip_22_27,ip_22_28,ip_22_29,ip_22_30,ip_22_31,ip_23_0,ip_23_1,ip_23_2,ip_23_3,ip_23_4,ip_23_5,ip_23_6,ip_23_7,ip_23_8,ip_23_9,ip_23_10,ip_23_11,ip_23_12,ip_23_13,ip_23_14,ip_23_15,ip_23_16,ip_23_17,ip_23_18,ip_23_19,ip_23_20,ip_23_21,ip_23_22,ip_23_23,ip_23_24,ip_23_25,ip_23_26,ip_23_27,ip_23_28,ip_23_29,ip_23_30,ip_23_31,ip_24_0,ip_24_1,ip_24_2,ip_24_3,ip_24_4,ip_24_5,ip_24_6,ip_24_7,ip_24_8,ip_24_9,ip_24_10,ip_24_11,ip_24_12,ip_24_13,ip_24_14,ip_24_15,ip_24_16,ip_24_17,ip_24_18,ip_24_19,ip_24_20,ip_24_21,ip_24_22,ip_24_23,ip_24_24,ip_24_25,ip_24_26,ip_24_27,ip_24_28,ip_24_29,ip_24_30,ip_24_31,ip_25_0,ip_25_1,ip_25_2,ip_25_3,ip_25_4,ip_25_5,ip_25_6,ip_25_7,ip_25_8,ip_25_9,ip_25_10,ip_25_11,ip_25_12,ip_25_13,ip_25_14,ip_25_15,ip_25_16,ip_25_17,ip_25_18,ip_25_19,ip_25_20,ip_25_21,ip_25_22,ip_25_23,ip_25_24,ip_25_25,ip_25_26,ip_25_27,ip_25_28,ip_25_29,ip_25_30,ip_25_31,ip_26_0,ip_26_1,ip_26_2,ip_26_3,ip_26_4,ip_26_5,ip_26_6,ip_26_7,ip_26_8,ip_26_9,ip_26_10,ip_26_11,ip_26_12,ip_26_13,ip_26_14,ip_26_15,ip_26_16,ip_26_17,ip_26_18,ip_26_19,ip_26_20,ip_26_21,ip_26_22,ip_26_23,ip_26_24,ip_26_25,ip_26_26,ip_26_27,ip_26_28,ip_26_29,ip_26_30,ip_26_31,ip_27_0,ip_27_1,ip_27_2,ip_27_3,ip_27_4,ip_27_5,ip_27_6,ip_27_7,ip_27_8,ip_27_9,ip_27_10,ip_27_11,ip_27_12,ip_27_13,ip_27_14,ip_27_15,ip_27_16,ip_27_17,ip_27_18,ip_27_19,ip_27_20,ip_27_21,ip_27_22,ip_27_23,ip_27_24,ip_27_25,ip_27_26,ip_27_27,ip_27_28,ip_27_29,ip_27_30,ip_27_31,ip_28_0,ip_28_1,ip_28_2,ip_28_3,ip_28_4,ip_28_5,ip_28_6,ip_28_7,ip_28_8,ip_28_9,ip_28_10,ip_28_11,ip_28_12,ip_28_13,ip_28_14,ip_28_15,ip_28_16,ip_28_17,ip_28_18,ip_28_19,ip_28_20,ip_28_21,ip_28_22,ip_28_23,ip_28_24,ip_28_25,ip_28_26,ip_28_27,ip_28_28,ip_28_29,ip_28_30,ip_28_31,ip_29_0,ip_29_1,ip_29_2,ip_29_3,ip_29_4,ip_29_5,ip_29_6,ip_29_7,ip_29_8,ip_29_9,ip_29_10,ip_29_11,ip_29_12,ip_29_13,ip_29_14,ip_29_15,ip_29_16,ip_29_17,ip_29_18,ip_29_19,ip_29_20,ip_29_21,ip_29_22,ip_29_23,ip_29_24,ip_29_25,ip_29_26,ip_29_27,ip_29_28,ip_29_29,ip_29_30,ip_29_31,ip_30_0,ip_30_1,ip_30_2,ip_30_3,ip_30_4,ip_30_5,ip_30_6,ip_30_7,ip_30_8,ip_30_9,ip_30_10,ip_30_11,ip_30_12,ip_30_13,ip_30_14,ip_30_15,ip_30_16,ip_30_17,ip_30_18,ip_30_19,ip_30_20,ip_30_21,ip_30_22,ip_30_23,ip_30_24,ip_30_25,ip_30_26,ip_30_27,ip_30_28,ip_30_29,ip_30_30,ip_30_31,ip_31_0,ip_31_1,ip_31_2,ip_31_3,ip_31_4,ip_31_5,ip_31_6,ip_31_7,ip_31_8,ip_31_9,ip_31_10,ip_31_11,ip_31_12,ip_31_13,ip_31_14,ip_31_15,ip_31_16,ip_31_17,ip_31_18,ip_31_19,ip_31_20,ip_31_21,ip_31_22,ip_31_23,ip_31_24,ip_31_25,ip_31_26,ip_31_27,ip_31_28,ip_31_29,ip_31_30,ip_31_31;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149,p1150,p1151,p1152,p1153,p1154,p1155,p1156,p1157,p1158,p1159,p1160,p1161,p1162,p1163,p1164,p1165,p1166,p1167,p1168,p1169,p1170,p1171,p1172,p1173,p1174,p1175,p1176,p1177,p1178,p1179,p1180,p1181,p1182,p1183,p1184,p1185,p1186,p1187,p1188,p1189,p1190,p1191,p1192,p1193,p1194,p1195,p1196,p1197,p1198,p1199,p1200,p1201,p1202,p1203,p1204,p1205,p1206,p1207,p1208,p1209,p1210,p1211,p1212,p1213,p1214,p1215,p1216,p1217,p1218,p1219,p1220,p1221,p1222,p1223,p1224,p1225,p1226,p1227,p1228,p1229,p1230,p1231,p1232,p1233,p1234,p1235,p1236,p1237,p1238,p1239,p1240,p1241,p1242,p1243,p1244,p1245,p1246,p1247,p1248,p1249,p1250,p1251,p1252,p1253,p1254,p1255,p1256,p1257,p1258,p1259,p1260,p1261,p1262,p1263,p1264,p1265,p1266,p1267,p1268,p1269,p1270,p1271,p1272,p1273,p1274,p1275,p1276,p1277,p1278,p1279,p1280,p1281,p1282,p1283,p1284,p1285,p1286,p1287,p1288,p1289,p1290,p1291,p1292,p1293,p1294,p1295,p1296,p1297,p1298,p1299,p1300,p1301,p1302,p1303,p1304,p1305,p1306,p1307,p1308,p1309,p1310,p1311,p1312,p1313,p1314,p1315,p1316,p1317,p1318,p1319,p1320,p1321,p1322,p1323,p1324,p1325,p1326,p1327,p1328,p1329,p1330,p1331,p1332,p1333,p1334,p1335,p1336,p1337,p1338,p1339,p1340,p1341,p1342,p1343,p1344,p1345,p1346,p1347,p1348,p1349,p1350,p1351,p1352,p1353,p1354,p1355,p1356,p1357,p1358,p1359,p1360,p1361,p1362,p1363,p1364,p1365,p1366,p1367,p1368,p1369,p1370,p1371,p1372,p1373,p1374,p1375,p1376,p1377,p1378,p1379,p1380,p1381,p1382,p1383,p1384,p1385,p1386,p1387,p1388,p1389,p1390,p1391,p1392,p1393,p1394,p1395,p1396,p1397,p1398,p1399,p1400,p1401,p1402,p1403,p1404,p1405,p1406,p1407,p1408,p1409,p1410,p1411,p1412,p1413,p1414,p1415,p1416,p1417,p1418,p1419,p1420,p1421,p1422,p1423,p1424,p1425,p1426,p1427,p1428,p1429,p1430,p1431,p1432,p1433,p1434,p1435,p1436,p1437,p1438,p1439,p1440,p1441,p1442,p1443,p1444,p1445,p1446,p1447,p1448,p1449,p1450,p1451,p1452,p1453,p1454,p1455,p1456,p1457,p1458,p1459,p1460,p1461,p1462,p1463,p1464,p1465,p1466,p1467,p1468,p1469,p1470,p1471,p1472,p1473,p1474,p1475,p1476,p1477,p1478,p1479,p1480,p1481,p1482,p1483,p1484,p1485,p1486,p1487,p1488,p1489,p1490,p1491,p1492,p1493,p1494,p1495,p1496,p1497,p1498,p1499,p1500,p1501,p1502,p1503,p1504,p1505,p1506,p1507,p1508,p1509,p1510,p1511,p1512,p1513,p1514,p1515,p1516,p1517,p1518,p1519,p1520,p1521,p1522,p1523,p1524,p1525,p1526,p1527,p1528,p1529,p1530,p1531,p1532,p1533,p1534,p1535,p1536,p1537,p1538,p1539,p1540,p1541,p1542,p1543,p1544,p1545,p1546,p1547,p1548,p1549,p1550,p1551,p1552,p1553,p1554,p1555,p1556,p1557,p1558,p1559,p1560,p1561,p1562,p1563,p1564,p1565,p1566,p1567,p1568,p1569,p1570,p1571,p1572,p1573,p1574,p1575,p1576,p1577,p1578,p1579,p1580,p1581,p1582,p1583,p1584,p1585,p1586,p1587,p1588,p1589,p1590,p1591,p1592,p1593,p1594,p1595,p1596,p1597,p1598,p1599,p1600,p1601,p1602,p1603,p1604,p1605,p1606,p1607,p1608,p1609,p1610,p1611,p1612,p1613,p1614,p1615,p1616,p1617,p1618,p1619,p1620,p1621,p1622,p1623,p1624,p1625,p1626,p1627,p1628,p1629,p1630,p1631,p1632,p1633,p1634,p1635,p1636,p1637,p1638,p1639,p1640,p1641,p1642,p1643,p1644,p1645,p1646,p1647,p1648,p1649,p1650,p1651,p1652,p1653,p1654,p1655,p1656,p1657,p1658,p1659,p1660,p1661,p1662,p1663,p1664,p1665,p1666,p1667,p1668,p1669,p1670,p1671,p1672,p1673,p1674,p1675,p1676,p1677,p1678,p1679,p1680,p1681,p1682,p1683,p1684,p1685,p1686,p1687,p1688,p1689,p1690,p1691,p1692,p1693,p1694,p1695,p1696,p1697,p1698,p1699,p1700,p1701,p1702,p1703,p1704,p1705,p1706,p1707,p1708,p1709,p1710,p1711,p1712,p1713,p1714,p1715,p1716,p1717,p1718,p1719,p1720,p1721,p1722,p1723,p1724,p1725,p1726,p1727,p1728,p1729,p1730,p1731,p1732,p1733,p1734,p1735,p1736,p1737,p1738,p1739,p1740,p1741,p1742,p1743,p1744,p1745,p1746,p1747,p1748,p1749,p1750,p1751,p1752,p1753,p1754,p1755,p1756,p1757,p1758,p1759,p1760,p1761,p1762,p1763,p1764,p1765,p1766,p1767,p1768,p1769,p1770,p1771,p1772,p1773,p1774,p1775,p1776,p1777,p1778,p1779,p1780,p1781,p1782,p1783,p1784,p1785,p1786,p1787,p1788,p1789,p1790,p1791,p1792,p1793,p1794,p1795,p1796,p1797,p1798,p1799,p1800,p1801,p1802,p1803,p1804,p1805,p1806,p1807,p1808,p1809,p1810,p1811,p1812,p1813,p1814,p1815,p1816,p1817,p1818,p1819,p1820,p1821,p1822,p1823,p1824,p1825,p1826,p1827,p1828,p1829,p1830,p1831,p1832,p1833,p1834,p1835,p1836,p1837,p1838,p1839,p1840,p1841,p1842,p1843,p1844,p1845,p1846,p1847,p1848,p1849,p1850,p1851,p1852,p1853,p1854,p1855,p1856,p1857,p1858,p1859,p1860,p1861,p1862,p1863,p1864,p1865,p1866,p1867,p1868,p1869,p1870,p1871,p1872,p1873,p1874,p1875,p1876,p1877,p1878,p1879,p1880,p1881,p1882,p1883,p1884,p1885,p1886,p1887,p1888,p1889,p1890,p1891,p1892,p1893,p1894,p1895,p1896,p1897,p1898,p1899,p1900,p1901,p1902,p1903,p1904,p1905,p1906,p1907,p1908,p1909,p1910,p1911,p1912,p1913,p1914,p1915,p1916,p1917,p1918,p1919,p1920,p1921,p1922,p1923,p1924,p1925,p1926,p1927,p1928,p1929,p1930,p1931,p1932,p1933,p1934,p1935,p1936,p1937,p1938,p1939,p1940,p1941,p1942,p1943,p1944,p1945,p1946,p1947,p1948,p1949,p1950,p1951,p1952,p1953,p1954,p1955,p1956,p1957,p1958,p1959,p1960,p1961,p1962,p1963,p1964,p1965,p1966,p1967,p1968,p1969,p1970,p1971,p1972,p1973,p1974,p1975,p1976,p1977,p1978,p1979,p1980,p1981,p1982,p1983,p1984,p1985,p1986,p1987,p1988,p1989,p1990,p1991,p1992,p1993,p1994,p1995,p1996,p1997,p1998,p1999,p2000,p2001,p2002,p2003,p2004,p2005,p2006,p2007,p2008,p2009,p2010,p2011,p2012,p2013,p2014,p2015,p2016,p2017,p2018,p2019,p2020,p2021,p2022,p2023,p2024,p2025,p2026,p2027,p2028,p2029,p2030,p2031,p2032,p2033,p2034,p2035,p2036,p2037,p2038,p2039,p2040,p2041,p2042,p2043,p2044,p2045,p2046,p2047,p2048,p2049,p2050,p2051,p2052,p2053,p2054,p2055,p2056,p2057,p2058,p2059,p2060,p2061,p2062,p2063,p2064,p2065,p2066,p2067,p2068,p2069,p2070,p2071,p2072,p2073,p2074,p2075,p2076,p2077,p2078,p2079,p2080,p2081,p2082,p2083,p2084,p2085,p2086,p2087,p2088,p2089,p2090,p2091,p2092,p2093,p2094,p2095,p2096,p2097,p2098,p2099,p2100,p2101,p2102,p2103,p2104,p2105,p2106,p2107,p2108,p2109,p2110,p2111,p2112,p2113,p2114,p2115,p2116,p2117,p2118,p2119,p2120,p2121,p2122,p2123,p2124,p2125,p2126,p2127,p2128,p2129,p2130,p2131,p2132,p2133,p2134,p2135,p2136,p2137,p2138,p2139,p2140,p2141,p2142,p2143,p2144,p2145,p2146,p2147,p2148,p2149,p2150,p2151,p2152,p2153,p2154,p2155,p2156,p2157,p2158,p2159,p2160,p2161,p2162,p2163,p2164,p2165,p2166,p2167,p2168,p2169,p2170,p2171,p2172,p2173,p2174,p2175,p2176,p2177,p2178,p2179,p2180,p2181,p2182,p2183,p2184,p2185,p2186,p2187,p2188,p2189,p2190,p2191,p2192,p2193,p2194,p2195,p2196,p2197,p2198,p2199,p2200,p2201,p2202,p2203,p2204,p2205,p2206,p2207,p2208,p2209,p2210,p2211,p2212,p2213,p2214,p2215,p2216,p2217,p2218,p2219,p2220,p2221,p2222,p2223,p2224,p2225,p2226,p2227,p2228,p2229,p2230,p2231,p2232,p2233,p2234,p2235,p2236,p2237,p2238,p2239,p2240,p2241,p2242,p2243,p2244,p2245,p2246,p2247,p2248,p2249,p2250,p2251,p2252,p2253,p2254,p2255,p2256,p2257,p2258,p2259,p2260,p2261,p2262,p2263,p2264,p2265,p2266,p2267,p2268,p2269,p2270,p2271,p2272,p2273,p2274,p2275,p2276,p2277,p2278,p2279,p2280,p2281,p2282,p2283,p2284,p2285,p2286,p2287,p2288,p2289,p2290,p2291,p2292,p2293,p2294,p2295,p2296,p2297,p2298,p2299,p2300,p2301,p2302,p2303,p2304,p2305,p2306,p2307,p2308,p2309,p2310,p2311,p2312,p2313,p2314,p2315,p2316,p2317,p2318,p2319,p2320,p2321,p2322,p2323,p2324,p2325,p2326,p2327,p2328,p2329,p2330,p2331,p2332,p2333,p2334,p2335,p2336,p2337,p2338,p2339,p2340,p2341,p2342,p2343,p2344,p2345,p2346,p2347,p2348,p2349,p2350,p2351,p2352,p2353,p2354,p2355,p2356,p2357,p2358,p2359,p2360,p2361,p2362,p2363,p2364,p2365,p2366,p2367,p2368,p2369,p2370,p2371,p2372,p2373,p2374,p2375,p2376,p2377,p2378,p2379,p2380,p2381,p2382,p2383,p2384,p2385,p2386,p2387,p2388,p2389,p2390,p2391,p2392,p2393,p2394,p2395,p2396,p2397,p2398,p2399,p2400,p2401,p2402,p2403,p2404,p2405,p2406,p2407,p2408,p2409,p2410,p2411,p2412,p2413,p2414,p2415,p2416,p2417,p2418,p2419,p2420,p2421,p2422,p2423,p2424,p2425,p2426,p2427,p2428,p2429,p2430,p2431,p2432,p2433,p2434,p2435,p2436,p2437,p2438,p2439,p2440,p2441,p2442,p2443,p2444,p2445,p2446,p2447,p2448,p2449,p2450,p2451,p2452,p2453,p2454,p2455,p2456,p2457,p2458,p2459,p2460,p2461,p2462,p2463,p2464,p2465,p2466,p2467,p2468,p2469,p2470,p2471,p2472,p2473,p2474,p2475,p2476,p2477,p2478,p2479,p2480,p2481,p2482,p2483,p2484,p2485,p2486,p2487,p2488,p2489,p2490,p2491,p2492,p2493,p2494,p2495,p2496,p2497,p2498,p2499,p2500,p2501,p2502,p2503,p2504,p2505,p2506,p2507,p2508,p2509,p2510,p2511,p2512,p2513,p2514,p2515,p2516,p2517,p2518,p2519,p2520,p2521,p2522,p2523,p2524,p2525,p2526,p2527,p2528,p2529,p2530,p2531,p2532,p2533,p2534,p2535,p2536,p2537,p2538,p2539,p2540,p2541,p2542,p2543,p2544,p2545,p2546,p2547,p2548,p2549,p2550,p2551,p2552,p2553,p2554,p2555,p2556,p2557,p2558,p2559,p2560,p2561,p2562,p2563,p2564,p2565,p2566,p2567,p2568,p2569,p2570,p2571,p2572,p2573,p2574,p2575,p2576,p2577,p2578,p2579,p2580,p2581,p2582,p2583,p2584,p2585,p2586,p2587,p2588,p2589,p2590,p2591,p2592,p2593,p2594,p2595,p2596,p2597,p2598,p2599,p2600,p2601,p2602,p2603,p2604,p2605,p2606,p2607,p2608,p2609,p2610,p2611,p2612,p2613,p2614,p2615,p2616,p2617,p2618,p2619,p2620,p2621,p2622,p2623,p2624,p2625,p2626,p2627,p2628,p2629,p2630,p2631,p2632,p2633,p2634,p2635,p2636,p2637,p2638,p2639,p2640,p2641,p2642,p2643,p2644,p2645,p2646,p2647,p2648,p2649,p2650,p2651,p2652,p2653,p2654,p2655,p2656,p2657,p2658,p2659,p2660,p2661,p2662,p2663,p2664,p2665,p2666,p2667,p2668,p2669,p2670,p2671,p2672,p2673,p2674,p2675,p2676,p2677,p2678,p2679,p2680,p2681,p2682,p2683,p2684,p2685,p2686,p2687,p2688,p2689,p2690,p2691,p2692,p2693,p2694,p2695,p2696,p2697,p2698,p2699,p2700,p2701,p2702,p2703,p2704,p2705,p2706,p2707,p2708,p2709,p2710,p2711,p2712,p2713,p2714,p2715,p2716,p2717,p2718,p2719,p2720,p2721,p2722,p2723,p2724,p2725,p2726,p2727,p2728,p2729,p2730,p2731,p2732,p2733,p2734,p2735,p2736,p2737,p2738,p2739,p2740,p2741,p2742,p2743,p2744,p2745,p2746,p2747,p2748,p2749,p2750,p2751,p2752,p2753,p2754,p2755,p2756,p2757,p2758,p2759,p2760,p2761,p2762,p2763,p2764,p2765,p2766,p2767,p2768,p2769,p2770,p2771,p2772,p2773,p2774,p2775,p2776,p2777,p2778,p2779,p2780,p2781,p2782,p2783,p2784,p2785,p2786,p2787,p2788,p2789,p2790,p2791,p2792,p2793,p2794,p2795,p2796,p2797,p2798,p2799,p2800,p2801,p2802,p2803,p2804,p2805,p2806,p2807,p2808,p2809,p2810,p2811,p2812,p2813,p2814,p2815,p2816,p2817,p2818,p2819,p2820,p2821,p2822,p2823,p2824,p2825,p2826,p2827,p2828,p2829,p2830,p2831,p2832,p2833,p2834,p2835,p2836,p2837,p2838,p2839,p2840,p2841,p2842,p2843,p2844,p2845,p2846,p2847,p2848,p2849,p2850,p2851,p2852,p2853,p2854,p2855,p2856,p2857,p2858,p2859,p2860,p2861,p2862,p2863,p2864,p2865,p2866,p2867,p2868,p2869,p2870,p2871,p2872,p2873,p2874,p2875,p2876,p2877,p2878,p2879,p2880,p2881,p2882,p2883,p2884,p2885,p2886,p2887,p2888,p2889,p2890,p2891,p2892,p2893,p2894,p2895,p2896,p2897,p2898,p2899,p2900,p2901,p2902,p2903,p2904,p2905,p2906,p2907,p2908,p2909,p2910,p2911,p2912,p2913,p2914,p2915,p2916,p2917,p2918,p2919,p2920,p2921,p2922,p2923,p2924,p2925,p2926,p2927,p2928,p2929,p2930,p2931,p2932,p2933,p2934,p2935,p2936,p2937,p2938,p2939,p2940,p2941,p2942,p2943,p2944,p2945,p2946,p2947,p2948,p2949,p2950,p2951,p2952,p2953,p2954,p2955,p2956,p2957,p2958,p2959,p2960,p2961,p2962,p2963,p2964,p2965,p2966,p2967,p2968,p2969,p2970,p2971,p2972,p2973,p2974,p2975,p2976,p2977,p2978,p2979,p2980,p2981,p2982,p2983,p2984,p2985,p2986,p2987,p2988,p2989,p2990,p2991,p2992,p2993,p2994,p2995,p2996,p2997,p2998,p2999,p3000,p3001,p3002,p3003,p3004,p3005,p3006,p3007,p3008,p3009,p3010,p3011,p3012,p3013,p3014,p3015,p3016,p3017,p3018,p3019,p3020,p3021,p3022,p3023,p3024,p3025,p3026,p3027,p3028,p3029,p3030,p3031,p3032,p3033,p3034,p3035,p3036,p3037,p3038,p3039,p3040,p3041,p3042,p3043,p3044,p3045,p3046,p3047,p3048,p3049,p3050,p3051,p3052,p3053,p3054,p3055,p3056,p3057,p3058,p3059,p3060,p3061,p3062,p3063,p3064,p3065,p3066,p3067,p3068,p3069,p3070,p3071,p3072,p3073,p3074,p3075,p3076,p3077,p3078,p3079,p3080,p3081,p3082,p3083,p3084,p3085,p3086,p3087,p3088,p3089,p3090,p3091,p3092,p3093,p3094,p3095,p3096,p3097,p3098,p3099,p3100,p3101,p3102,p3103,p3104,p3105,p3106,p3107,p3108,p3109,p3110,p3111,p3112,p3113,p3114,p3115,p3116,p3117,p3118,p3119,p3120,p3121,p3122,p3123,p3124,p3125,p3126,p3127,p3128,p3129,p3130,p3131,p3132,p3133,p3134,p3135,p3136,p3137,p3138,p3139,p3140,p3141,p3142,p3143,p3144,p3145,p3146,p3147,p3148,p3149,p3150,p3151,p3152,p3153,p3154,p3155,p3156,p3157,p3158,p3159,p3160,p3161,p3162,p3163,p3164,p3165,p3166,p3167,p3168,p3169,p3170,p3171,p3172,p3173,p3174,p3175,p3176,p3177,p3178,p3179,p3180,p3181,p3182,p3183,p3184,p3185,p3186,p3187,p3188,p3189,p3190,p3191,p3192,p3193,p3194,p3195,p3196,p3197,p3198,p3199,p3200,p3201,p3202,p3203,p3204,p3205,p3206,p3207,p3208,p3209,p3210,p3211,p3212,p3213,p3214,p3215,p3216,p3217,p3218,p3219,p3220,p3221,p3222,p3223,p3224,p3225,p3226,p3227,p3228,p3229,p3230,p3231,p3232,p3233,p3234,p3235,p3236,p3237,p3238,p3239,p3240,p3241,p3242,p3243,p3244,p3245,p3246,p3247,p3248,p3249,p3250,p3251,p3252,p3253,p3254,p3255,p3256,p3257,p3258,p3259,p3260,p3261,p3262,p3263,p3264,p3265,p3266,p3267,p3268,p3269,p3270,p3271,p3272,p3273,p3274,p3275,p3276,p3277,p3278,p3279,p3280,p3281,p3282,p3283,p3284,p3285,p3286,p3287,p3288,p3289,p3290,p3291,p3292,p3293,p3294,p3295,p3296,p3297,p3298,p3299,p3300,p3301,p3302,p3303,p3304,p3305,p3306,p3307,p3308,p3309,p3310,p3311,p3312,p3313,p3314,p3315,p3316,p3317,p3318,p3319,p3320,p3321,p3322,p3323,p3324,p3325,p3326,p3327,p3328,p3329,p3330,p3331,p3332,p3333,p3334,p3335,p3336,p3337,p3338,p3339,p3340,p3341,p3342,p3343,p3344,p3345,p3346,p3347,p3348,p3349,p3350,p3351,p3352,p3353,p3354,p3355,p3356,p3357,p3358,p3359,p3360,p3361,p3362,p3363,p3364,p3365,p3366,p3367,p3368,p3369,p3370,p3371,p3372,p3373,p3374,p3375,p3376,p3377,p3378,p3379,p3380,p3381,p3382,p3383,p3384,p3385,p3386,p3387,p3388,p3389,p3390,p3391,p3392,p3393,p3394,p3395,p3396,p3397,p3398,p3399,p3400,p3401,p3402,p3403,p3404,p3405,p3406,p3407,p3408,p3409,p3410,p3411,p3412,p3413,p3414,p3415,p3416,p3417,p3418,p3419,p3420,p3421,p3422,p3423,p3424,p3425,p3426,p3427,p3428,p3429,p3430,p3431,p3432,p3433,p3434,p3435,p3436,p3437,p3438,p3439,p3440,p3441,p3442,p3443,p3444,p3445,p3446,p3447,p3448,p3449,p3450,p3451,p3452,p3453,p3454,p3455,p3456,p3457,p3458,p3459,p3460,p3461,p3462,p3463,p3464,p3465,p3466,p3467,p3468,p3469,p3470,p3471,p3472,p3473,p3474,p3475,p3476,p3477,p3478,p3479,p3480,p3481,p3482,p3483,p3484,p3485,p3486,p3487,p3488,p3489,p3490,p3491,p3492,p3493,p3494,p3495,p3496,p3497,p3498,p3499,p3500,p3501,p3502,p3503,p3504,p3505,p3506,p3507,p3508,p3509,p3510,p3511,p3512,p3513,p3514,p3515,p3516,p3517,p3518,p3519,p3520,p3521,p3522,p3523,p3524,p3525,p3526,p3527,p3528,p3529,p3530,p3531,p3532,p3533,p3534,p3535,p3536,p3537,p3538,p3539,p3540,p3541,p3542,p3543,p3544,p3545,p3546,p3547,p3548,p3549,p3550,p3551,p3552,p3553,p3554,p3555,p3556,p3557,p3558,p3559,p3560,p3561,p3562,p3563,p3564,p3565,p3566,p3567,p3568,p3569,p3570,p3571,p3572,p3573,p3574,p3575,p3576,p3577,p3578,p3579,p3580,p3581,p3582,p3583,p3584,p3585,p3586,p3587,p3588,p3589,p3590,p3591,p3592,p3593,p3594,p3595,p3596,p3597,p3598,p3599,p3600,p3601,p3602,p3603,p3604,p3605,p3606,p3607,p3608,p3609,p3610,p3611,p3612,p3613,p3614,p3615,p3616,p3617,p3618,p3619,p3620,p3621,p3622,p3623,p3624,p3625,p3626,p3627,p3628,p3629,p3630,p3631,p3632,p3633,p3634,p3635,p3636,p3637,p3638,p3639,p3640,p3641,p3642,p3643,p3644,p3645,p3646,p3647,p3648,p3649,p3650,p3651,p3652,p3653,p3654,p3655,p3656,p3657,p3658,p3659,p3660,p3661,p3662,p3663,p3664,p3665,p3666,p3667,p3668,p3669,p3670,p3671,p3672,p3673,p3674,p3675,p3676,p3677,p3678,p3679,p3680,p3681,p3682,p3683,p3684,p3685,p3686,p3687,p3688,p3689,p3690,p3691,p3692,p3693,p3694,p3695,p3696,p3697,p3698,p3699,p3700,p3701,p3702,p3703,p3704,p3705,p3706,p3707,p3708,p3709,p3710,p3711,p3712,p3713,p3714,p3715,p3716,p3717,p3718,p3719,p3720,p3721,p3722,p3723,p3724,p3725,p3726,p3727,p3728,p3729,p3730,p3731,p3732,p3733,p3734,p3735,p3736,p3737,p3738,p3739,p3740,p3741,p3742,p3743,p3744,p3745,p3746,p3747,p3748,p3749,p3750,p3751,p3752,p3753,p3754,p3755,p3756,p3757,p3758,p3759,p3760,p3761,p3762,p3763,p3764,p3765,p3766,p3767,p3768,p3769,p3770,p3771,p3772,p3773,p3774,p3775,p3776,p3777,p3778,p3779,p3780,p3781,p3782,p3783,p3784,p3785,p3786,p3787,p3788,p3789,p3790,p3791,p3792,p3793,p3794,p3795,p3796,p3797,p3798,p3799,p3800,p3801,p3802,p3803,p3804,p3805,p3806,p3807,p3808,p3809,p3810,p3811,p3812,p3813,p3814,p3815,p3816,p3817,p3818,p3819,p3820,p3821,p3822,p3823,p3824,p3825,p3826,p3827,p3828,p3829,p3830,p3831,p3832,p3833,p3834,p3835,p3836,p3837,p3838,p3839,p3840,p3841,p3842,p3843,p3844,p3845,p3846,p3847,p3848,p3849,p3850,p3851,p3852,p3853,p3854,p3855,p3856,p3857,p3858,p3859,p3860,p3861,p3862,p3863,p3864,p3865,p3866,p3867,p3868,p3869,p3870,p3871,p3872,p3873,p3874,p3875,p3876,p3877,p3878,p3879,p3880,p3881,p3882,p3883,p3884,p3885,p3886,p3887,p3888,p3889,p3890,p3891,p3892,p3893,p3894,p3895,p3896,p3897,p3898,p3899,p3900,p3901,p3902,p3903,p3904,p3905,p3906,p3907,p3908,p3909,p3910,p3911,p3912,p3913,p3914,p3915,p3916,p3917,p3918,p3919,p3920,p3921,p3922,p3923,p3924,p3925,p3926,p3927,p3928,p3929,p3930,p3931,p3932,p3933,p3934,p3935,p3936,p3937,p3938,p3939,p3940,p3941,p3942,p3943,p3944,p3945,p3946,p3947,p3948,p3949,p3950,p3951,p3952,p3953,p3954,p3955,p3956,p3957,p3958,p3959,p3960,p3961,p3962,p3963,p3964,p3965,p3966,p3967,p3968,p3969,p3970,p3971,p3972,p3973,p3974,p3975,p3976,p3977;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_0_16,x[0],y[16]);
and and17(ip_0_17,x[0],y[17]);
and and18(ip_0_18,x[0],y[18]);
and and19(ip_0_19,x[0],y[19]);
and and20(ip_0_20,x[0],y[20]);
and and21(ip_0_21,x[0],y[21]);
and and22(ip_0_22,x[0],y[22]);
and and23(ip_0_23,x[0],y[23]);
and and24(ip_0_24,x[0],y[24]);
and and25(ip_0_25,x[0],y[25]);
and and26(ip_0_26,x[0],y[26]);
and and27(ip_0_27,x[0],y[27]);
and and28(ip_0_28,x[0],y[28]);
and and29(ip_0_29,x[0],y[29]);
and and30(ip_0_30,x[0],y[30]);
and and31(ip_0_31,x[0],y[31]);
and and32(ip_1_0,x[1],y[0]);
and and33(ip_1_1,x[1],y[1]);
and and34(ip_1_2,x[1],y[2]);
and and35(ip_1_3,x[1],y[3]);
and and36(ip_1_4,x[1],y[4]);
and and37(ip_1_5,x[1],y[5]);
and and38(ip_1_6,x[1],y[6]);
and and39(ip_1_7,x[1],y[7]);
and and40(ip_1_8,x[1],y[8]);
and and41(ip_1_9,x[1],y[9]);
and and42(ip_1_10,x[1],y[10]);
and and43(ip_1_11,x[1],y[11]);
and and44(ip_1_12,x[1],y[12]);
and and45(ip_1_13,x[1],y[13]);
and and46(ip_1_14,x[1],y[14]);
and and47(ip_1_15,x[1],y[15]);
and and48(ip_1_16,x[1],y[16]);
and and49(ip_1_17,x[1],y[17]);
and and50(ip_1_18,x[1],y[18]);
and and51(ip_1_19,x[1],y[19]);
and and52(ip_1_20,x[1],y[20]);
and and53(ip_1_21,x[1],y[21]);
and and54(ip_1_22,x[1],y[22]);
and and55(ip_1_23,x[1],y[23]);
and and56(ip_1_24,x[1],y[24]);
and and57(ip_1_25,x[1],y[25]);
and and58(ip_1_26,x[1],y[26]);
and and59(ip_1_27,x[1],y[27]);
and and60(ip_1_28,x[1],y[28]);
and and61(ip_1_29,x[1],y[29]);
and and62(ip_1_30,x[1],y[30]);
and and63(ip_1_31,x[1],y[31]);
and and64(ip_2_0,x[2],y[0]);
and and65(ip_2_1,x[2],y[1]);
and and66(ip_2_2,x[2],y[2]);
and and67(ip_2_3,x[2],y[3]);
and and68(ip_2_4,x[2],y[4]);
and and69(ip_2_5,x[2],y[5]);
and and70(ip_2_6,x[2],y[6]);
and and71(ip_2_7,x[2],y[7]);
and and72(ip_2_8,x[2],y[8]);
and and73(ip_2_9,x[2],y[9]);
and and74(ip_2_10,x[2],y[10]);
and and75(ip_2_11,x[2],y[11]);
and and76(ip_2_12,x[2],y[12]);
and and77(ip_2_13,x[2],y[13]);
and and78(ip_2_14,x[2],y[14]);
and and79(ip_2_15,x[2],y[15]);
and and80(ip_2_16,x[2],y[16]);
and and81(ip_2_17,x[2],y[17]);
and and82(ip_2_18,x[2],y[18]);
and and83(ip_2_19,x[2],y[19]);
and and84(ip_2_20,x[2],y[20]);
and and85(ip_2_21,x[2],y[21]);
and and86(ip_2_22,x[2],y[22]);
and and87(ip_2_23,x[2],y[23]);
and and88(ip_2_24,x[2],y[24]);
and and89(ip_2_25,x[2],y[25]);
and and90(ip_2_26,x[2],y[26]);
and and91(ip_2_27,x[2],y[27]);
and and92(ip_2_28,x[2],y[28]);
and and93(ip_2_29,x[2],y[29]);
and and94(ip_2_30,x[2],y[30]);
and and95(ip_2_31,x[2],y[31]);
and and96(ip_3_0,x[3],y[0]);
and and97(ip_3_1,x[3],y[1]);
and and98(ip_3_2,x[3],y[2]);
and and99(ip_3_3,x[3],y[3]);
and and100(ip_3_4,x[3],y[4]);
and and101(ip_3_5,x[3],y[5]);
and and102(ip_3_6,x[3],y[6]);
and and103(ip_3_7,x[3],y[7]);
and and104(ip_3_8,x[3],y[8]);
and and105(ip_3_9,x[3],y[9]);
and and106(ip_3_10,x[3],y[10]);
and and107(ip_3_11,x[3],y[11]);
and and108(ip_3_12,x[3],y[12]);
and and109(ip_3_13,x[3],y[13]);
and and110(ip_3_14,x[3],y[14]);
and and111(ip_3_15,x[3],y[15]);
and and112(ip_3_16,x[3],y[16]);
and and113(ip_3_17,x[3],y[17]);
and and114(ip_3_18,x[3],y[18]);
and and115(ip_3_19,x[3],y[19]);
and and116(ip_3_20,x[3],y[20]);
and and117(ip_3_21,x[3],y[21]);
and and118(ip_3_22,x[3],y[22]);
and and119(ip_3_23,x[3],y[23]);
and and120(ip_3_24,x[3],y[24]);
and and121(ip_3_25,x[3],y[25]);
and and122(ip_3_26,x[3],y[26]);
and and123(ip_3_27,x[3],y[27]);
and and124(ip_3_28,x[3],y[28]);
and and125(ip_3_29,x[3],y[29]);
and and126(ip_3_30,x[3],y[30]);
and and127(ip_3_31,x[3],y[31]);
and and128(ip_4_0,x[4],y[0]);
and and129(ip_4_1,x[4],y[1]);
and and130(ip_4_2,x[4],y[2]);
and and131(ip_4_3,x[4],y[3]);
and and132(ip_4_4,x[4],y[4]);
and and133(ip_4_5,x[4],y[5]);
and and134(ip_4_6,x[4],y[6]);
and and135(ip_4_7,x[4],y[7]);
and and136(ip_4_8,x[4],y[8]);
and and137(ip_4_9,x[4],y[9]);
and and138(ip_4_10,x[4],y[10]);
and and139(ip_4_11,x[4],y[11]);
and and140(ip_4_12,x[4],y[12]);
and and141(ip_4_13,x[4],y[13]);
and and142(ip_4_14,x[4],y[14]);
and and143(ip_4_15,x[4],y[15]);
and and144(ip_4_16,x[4],y[16]);
and and145(ip_4_17,x[4],y[17]);
and and146(ip_4_18,x[4],y[18]);
and and147(ip_4_19,x[4],y[19]);
and and148(ip_4_20,x[4],y[20]);
and and149(ip_4_21,x[4],y[21]);
and and150(ip_4_22,x[4],y[22]);
and and151(ip_4_23,x[4],y[23]);
and and152(ip_4_24,x[4],y[24]);
and and153(ip_4_25,x[4],y[25]);
and and154(ip_4_26,x[4],y[26]);
and and155(ip_4_27,x[4],y[27]);
and and156(ip_4_28,x[4],y[28]);
and and157(ip_4_29,x[4],y[29]);
and and158(ip_4_30,x[4],y[30]);
and and159(ip_4_31,x[4],y[31]);
and and160(ip_5_0,x[5],y[0]);
and and161(ip_5_1,x[5],y[1]);
and and162(ip_5_2,x[5],y[2]);
and and163(ip_5_3,x[5],y[3]);
and and164(ip_5_4,x[5],y[4]);
and and165(ip_5_5,x[5],y[5]);
and and166(ip_5_6,x[5],y[6]);
and and167(ip_5_7,x[5],y[7]);
and and168(ip_5_8,x[5],y[8]);
and and169(ip_5_9,x[5],y[9]);
and and170(ip_5_10,x[5],y[10]);
and and171(ip_5_11,x[5],y[11]);
and and172(ip_5_12,x[5],y[12]);
and and173(ip_5_13,x[5],y[13]);
and and174(ip_5_14,x[5],y[14]);
and and175(ip_5_15,x[5],y[15]);
and and176(ip_5_16,x[5],y[16]);
and and177(ip_5_17,x[5],y[17]);
and and178(ip_5_18,x[5],y[18]);
and and179(ip_5_19,x[5],y[19]);
and and180(ip_5_20,x[5],y[20]);
and and181(ip_5_21,x[5],y[21]);
and and182(ip_5_22,x[5],y[22]);
and and183(ip_5_23,x[5],y[23]);
and and184(ip_5_24,x[5],y[24]);
and and185(ip_5_25,x[5],y[25]);
and and186(ip_5_26,x[5],y[26]);
and and187(ip_5_27,x[5],y[27]);
and and188(ip_5_28,x[5],y[28]);
and and189(ip_5_29,x[5],y[29]);
and and190(ip_5_30,x[5],y[30]);
and and191(ip_5_31,x[5],y[31]);
and and192(ip_6_0,x[6],y[0]);
and and193(ip_6_1,x[6],y[1]);
and and194(ip_6_2,x[6],y[2]);
and and195(ip_6_3,x[6],y[3]);
and and196(ip_6_4,x[6],y[4]);
and and197(ip_6_5,x[6],y[5]);
and and198(ip_6_6,x[6],y[6]);
and and199(ip_6_7,x[6],y[7]);
and and200(ip_6_8,x[6],y[8]);
and and201(ip_6_9,x[6],y[9]);
and and202(ip_6_10,x[6],y[10]);
and and203(ip_6_11,x[6],y[11]);
and and204(ip_6_12,x[6],y[12]);
and and205(ip_6_13,x[6],y[13]);
and and206(ip_6_14,x[6],y[14]);
and and207(ip_6_15,x[6],y[15]);
and and208(ip_6_16,x[6],y[16]);
and and209(ip_6_17,x[6],y[17]);
and and210(ip_6_18,x[6],y[18]);
and and211(ip_6_19,x[6],y[19]);
and and212(ip_6_20,x[6],y[20]);
and and213(ip_6_21,x[6],y[21]);
and and214(ip_6_22,x[6],y[22]);
and and215(ip_6_23,x[6],y[23]);
and and216(ip_6_24,x[6],y[24]);
and and217(ip_6_25,x[6],y[25]);
and and218(ip_6_26,x[6],y[26]);
and and219(ip_6_27,x[6],y[27]);
and and220(ip_6_28,x[6],y[28]);
and and221(ip_6_29,x[6],y[29]);
and and222(ip_6_30,x[6],y[30]);
and and223(ip_6_31,x[6],y[31]);
and and224(ip_7_0,x[7],y[0]);
and and225(ip_7_1,x[7],y[1]);
and and226(ip_7_2,x[7],y[2]);
and and227(ip_7_3,x[7],y[3]);
and and228(ip_7_4,x[7],y[4]);
and and229(ip_7_5,x[7],y[5]);
and and230(ip_7_6,x[7],y[6]);
and and231(ip_7_7,x[7],y[7]);
and and232(ip_7_8,x[7],y[8]);
and and233(ip_7_9,x[7],y[9]);
and and234(ip_7_10,x[7],y[10]);
and and235(ip_7_11,x[7],y[11]);
and and236(ip_7_12,x[7],y[12]);
and and237(ip_7_13,x[7],y[13]);
and and238(ip_7_14,x[7],y[14]);
and and239(ip_7_15,x[7],y[15]);
and and240(ip_7_16,x[7],y[16]);
and and241(ip_7_17,x[7],y[17]);
and and242(ip_7_18,x[7],y[18]);
and and243(ip_7_19,x[7],y[19]);
and and244(ip_7_20,x[7],y[20]);
and and245(ip_7_21,x[7],y[21]);
and and246(ip_7_22,x[7],y[22]);
and and247(ip_7_23,x[7],y[23]);
and and248(ip_7_24,x[7],y[24]);
and and249(ip_7_25,x[7],y[25]);
and and250(ip_7_26,x[7],y[26]);
and and251(ip_7_27,x[7],y[27]);
and and252(ip_7_28,x[7],y[28]);
and and253(ip_7_29,x[7],y[29]);
and and254(ip_7_30,x[7],y[30]);
and and255(ip_7_31,x[7],y[31]);
and and256(ip_8_0,x[8],y[0]);
and and257(ip_8_1,x[8],y[1]);
and and258(ip_8_2,x[8],y[2]);
and and259(ip_8_3,x[8],y[3]);
and and260(ip_8_4,x[8],y[4]);
and and261(ip_8_5,x[8],y[5]);
and and262(ip_8_6,x[8],y[6]);
and and263(ip_8_7,x[8],y[7]);
and and264(ip_8_8,x[8],y[8]);
and and265(ip_8_9,x[8],y[9]);
and and266(ip_8_10,x[8],y[10]);
and and267(ip_8_11,x[8],y[11]);
and and268(ip_8_12,x[8],y[12]);
and and269(ip_8_13,x[8],y[13]);
and and270(ip_8_14,x[8],y[14]);
and and271(ip_8_15,x[8],y[15]);
and and272(ip_8_16,x[8],y[16]);
and and273(ip_8_17,x[8],y[17]);
and and274(ip_8_18,x[8],y[18]);
and and275(ip_8_19,x[8],y[19]);
and and276(ip_8_20,x[8],y[20]);
and and277(ip_8_21,x[8],y[21]);
and and278(ip_8_22,x[8],y[22]);
and and279(ip_8_23,x[8],y[23]);
and and280(ip_8_24,x[8],y[24]);
and and281(ip_8_25,x[8],y[25]);
and and282(ip_8_26,x[8],y[26]);
and and283(ip_8_27,x[8],y[27]);
and and284(ip_8_28,x[8],y[28]);
and and285(ip_8_29,x[8],y[29]);
and and286(ip_8_30,x[8],y[30]);
and and287(ip_8_31,x[8],y[31]);
and and288(ip_9_0,x[9],y[0]);
and and289(ip_9_1,x[9],y[1]);
and and290(ip_9_2,x[9],y[2]);
and and291(ip_9_3,x[9],y[3]);
and and292(ip_9_4,x[9],y[4]);
and and293(ip_9_5,x[9],y[5]);
and and294(ip_9_6,x[9],y[6]);
and and295(ip_9_7,x[9],y[7]);
and and296(ip_9_8,x[9],y[8]);
and and297(ip_9_9,x[9],y[9]);
and and298(ip_9_10,x[9],y[10]);
and and299(ip_9_11,x[9],y[11]);
and and300(ip_9_12,x[9],y[12]);
and and301(ip_9_13,x[9],y[13]);
and and302(ip_9_14,x[9],y[14]);
and and303(ip_9_15,x[9],y[15]);
and and304(ip_9_16,x[9],y[16]);
and and305(ip_9_17,x[9],y[17]);
and and306(ip_9_18,x[9],y[18]);
and and307(ip_9_19,x[9],y[19]);
and and308(ip_9_20,x[9],y[20]);
and and309(ip_9_21,x[9],y[21]);
and and310(ip_9_22,x[9],y[22]);
and and311(ip_9_23,x[9],y[23]);
and and312(ip_9_24,x[9],y[24]);
and and313(ip_9_25,x[9],y[25]);
and and314(ip_9_26,x[9],y[26]);
and and315(ip_9_27,x[9],y[27]);
and and316(ip_9_28,x[9],y[28]);
and and317(ip_9_29,x[9],y[29]);
and and318(ip_9_30,x[9],y[30]);
and and319(ip_9_31,x[9],y[31]);
and and320(ip_10_0,x[10],y[0]);
and and321(ip_10_1,x[10],y[1]);
and and322(ip_10_2,x[10],y[2]);
and and323(ip_10_3,x[10],y[3]);
and and324(ip_10_4,x[10],y[4]);
and and325(ip_10_5,x[10],y[5]);
and and326(ip_10_6,x[10],y[6]);
and and327(ip_10_7,x[10],y[7]);
and and328(ip_10_8,x[10],y[8]);
and and329(ip_10_9,x[10],y[9]);
and and330(ip_10_10,x[10],y[10]);
and and331(ip_10_11,x[10],y[11]);
and and332(ip_10_12,x[10],y[12]);
and and333(ip_10_13,x[10],y[13]);
and and334(ip_10_14,x[10],y[14]);
and and335(ip_10_15,x[10],y[15]);
and and336(ip_10_16,x[10],y[16]);
and and337(ip_10_17,x[10],y[17]);
and and338(ip_10_18,x[10],y[18]);
and and339(ip_10_19,x[10],y[19]);
and and340(ip_10_20,x[10],y[20]);
and and341(ip_10_21,x[10],y[21]);
and and342(ip_10_22,x[10],y[22]);
and and343(ip_10_23,x[10],y[23]);
and and344(ip_10_24,x[10],y[24]);
and and345(ip_10_25,x[10],y[25]);
and and346(ip_10_26,x[10],y[26]);
and and347(ip_10_27,x[10],y[27]);
and and348(ip_10_28,x[10],y[28]);
and and349(ip_10_29,x[10],y[29]);
and and350(ip_10_30,x[10],y[30]);
and and351(ip_10_31,x[10],y[31]);
and and352(ip_11_0,x[11],y[0]);
and and353(ip_11_1,x[11],y[1]);
and and354(ip_11_2,x[11],y[2]);
and and355(ip_11_3,x[11],y[3]);
and and356(ip_11_4,x[11],y[4]);
and and357(ip_11_5,x[11],y[5]);
and and358(ip_11_6,x[11],y[6]);
and and359(ip_11_7,x[11],y[7]);
and and360(ip_11_8,x[11],y[8]);
and and361(ip_11_9,x[11],y[9]);
and and362(ip_11_10,x[11],y[10]);
and and363(ip_11_11,x[11],y[11]);
and and364(ip_11_12,x[11],y[12]);
and and365(ip_11_13,x[11],y[13]);
and and366(ip_11_14,x[11],y[14]);
and and367(ip_11_15,x[11],y[15]);
and and368(ip_11_16,x[11],y[16]);
and and369(ip_11_17,x[11],y[17]);
and and370(ip_11_18,x[11],y[18]);
and and371(ip_11_19,x[11],y[19]);
and and372(ip_11_20,x[11],y[20]);
and and373(ip_11_21,x[11],y[21]);
and and374(ip_11_22,x[11],y[22]);
and and375(ip_11_23,x[11],y[23]);
and and376(ip_11_24,x[11],y[24]);
and and377(ip_11_25,x[11],y[25]);
and and378(ip_11_26,x[11],y[26]);
and and379(ip_11_27,x[11],y[27]);
and and380(ip_11_28,x[11],y[28]);
and and381(ip_11_29,x[11],y[29]);
and and382(ip_11_30,x[11],y[30]);
and and383(ip_11_31,x[11],y[31]);
and and384(ip_12_0,x[12],y[0]);
and and385(ip_12_1,x[12],y[1]);
and and386(ip_12_2,x[12],y[2]);
and and387(ip_12_3,x[12],y[3]);
and and388(ip_12_4,x[12],y[4]);
and and389(ip_12_5,x[12],y[5]);
and and390(ip_12_6,x[12],y[6]);
and and391(ip_12_7,x[12],y[7]);
and and392(ip_12_8,x[12],y[8]);
and and393(ip_12_9,x[12],y[9]);
and and394(ip_12_10,x[12],y[10]);
and and395(ip_12_11,x[12],y[11]);
and and396(ip_12_12,x[12],y[12]);
and and397(ip_12_13,x[12],y[13]);
and and398(ip_12_14,x[12],y[14]);
and and399(ip_12_15,x[12],y[15]);
and and400(ip_12_16,x[12],y[16]);
and and401(ip_12_17,x[12],y[17]);
and and402(ip_12_18,x[12],y[18]);
and and403(ip_12_19,x[12],y[19]);
and and404(ip_12_20,x[12],y[20]);
and and405(ip_12_21,x[12],y[21]);
and and406(ip_12_22,x[12],y[22]);
and and407(ip_12_23,x[12],y[23]);
and and408(ip_12_24,x[12],y[24]);
and and409(ip_12_25,x[12],y[25]);
and and410(ip_12_26,x[12],y[26]);
and and411(ip_12_27,x[12],y[27]);
and and412(ip_12_28,x[12],y[28]);
and and413(ip_12_29,x[12],y[29]);
and and414(ip_12_30,x[12],y[30]);
and and415(ip_12_31,x[12],y[31]);
and and416(ip_13_0,x[13],y[0]);
and and417(ip_13_1,x[13],y[1]);
and and418(ip_13_2,x[13],y[2]);
and and419(ip_13_3,x[13],y[3]);
and and420(ip_13_4,x[13],y[4]);
and and421(ip_13_5,x[13],y[5]);
and and422(ip_13_6,x[13],y[6]);
and and423(ip_13_7,x[13],y[7]);
and and424(ip_13_8,x[13],y[8]);
and and425(ip_13_9,x[13],y[9]);
and and426(ip_13_10,x[13],y[10]);
and and427(ip_13_11,x[13],y[11]);
and and428(ip_13_12,x[13],y[12]);
and and429(ip_13_13,x[13],y[13]);
and and430(ip_13_14,x[13],y[14]);
and and431(ip_13_15,x[13],y[15]);
and and432(ip_13_16,x[13],y[16]);
and and433(ip_13_17,x[13],y[17]);
and and434(ip_13_18,x[13],y[18]);
and and435(ip_13_19,x[13],y[19]);
and and436(ip_13_20,x[13],y[20]);
and and437(ip_13_21,x[13],y[21]);
and and438(ip_13_22,x[13],y[22]);
and and439(ip_13_23,x[13],y[23]);
and and440(ip_13_24,x[13],y[24]);
and and441(ip_13_25,x[13],y[25]);
and and442(ip_13_26,x[13],y[26]);
and and443(ip_13_27,x[13],y[27]);
and and444(ip_13_28,x[13],y[28]);
and and445(ip_13_29,x[13],y[29]);
and and446(ip_13_30,x[13],y[30]);
and and447(ip_13_31,x[13],y[31]);
and and448(ip_14_0,x[14],y[0]);
and and449(ip_14_1,x[14],y[1]);
and and450(ip_14_2,x[14],y[2]);
and and451(ip_14_3,x[14],y[3]);
and and452(ip_14_4,x[14],y[4]);
and and453(ip_14_5,x[14],y[5]);
and and454(ip_14_6,x[14],y[6]);
and and455(ip_14_7,x[14],y[7]);
and and456(ip_14_8,x[14],y[8]);
and and457(ip_14_9,x[14],y[9]);
and and458(ip_14_10,x[14],y[10]);
and and459(ip_14_11,x[14],y[11]);
and and460(ip_14_12,x[14],y[12]);
and and461(ip_14_13,x[14],y[13]);
and and462(ip_14_14,x[14],y[14]);
and and463(ip_14_15,x[14],y[15]);
and and464(ip_14_16,x[14],y[16]);
and and465(ip_14_17,x[14],y[17]);
and and466(ip_14_18,x[14],y[18]);
and and467(ip_14_19,x[14],y[19]);
and and468(ip_14_20,x[14],y[20]);
and and469(ip_14_21,x[14],y[21]);
and and470(ip_14_22,x[14],y[22]);
and and471(ip_14_23,x[14],y[23]);
and and472(ip_14_24,x[14],y[24]);
and and473(ip_14_25,x[14],y[25]);
and and474(ip_14_26,x[14],y[26]);
and and475(ip_14_27,x[14],y[27]);
and and476(ip_14_28,x[14],y[28]);
and and477(ip_14_29,x[14],y[29]);
and and478(ip_14_30,x[14],y[30]);
and and479(ip_14_31,x[14],y[31]);
and and480(ip_15_0,x[15],y[0]);
and and481(ip_15_1,x[15],y[1]);
and and482(ip_15_2,x[15],y[2]);
and and483(ip_15_3,x[15],y[3]);
and and484(ip_15_4,x[15],y[4]);
and and485(ip_15_5,x[15],y[5]);
and and486(ip_15_6,x[15],y[6]);
and and487(ip_15_7,x[15],y[7]);
and and488(ip_15_8,x[15],y[8]);
and and489(ip_15_9,x[15],y[9]);
and and490(ip_15_10,x[15],y[10]);
and and491(ip_15_11,x[15],y[11]);
and and492(ip_15_12,x[15],y[12]);
and and493(ip_15_13,x[15],y[13]);
and and494(ip_15_14,x[15],y[14]);
and and495(ip_15_15,x[15],y[15]);
and and496(ip_15_16,x[15],y[16]);
and and497(ip_15_17,x[15],y[17]);
and and498(ip_15_18,x[15],y[18]);
and and499(ip_15_19,x[15],y[19]);
and and500(ip_15_20,x[15],y[20]);
and and501(ip_15_21,x[15],y[21]);
and and502(ip_15_22,x[15],y[22]);
and and503(ip_15_23,x[15],y[23]);
and and504(ip_15_24,x[15],y[24]);
and and505(ip_15_25,x[15],y[25]);
and and506(ip_15_26,x[15],y[26]);
and and507(ip_15_27,x[15],y[27]);
and and508(ip_15_28,x[15],y[28]);
and and509(ip_15_29,x[15],y[29]);
and and510(ip_15_30,x[15],y[30]);
and and511(ip_15_31,x[15],y[31]);
and and512(ip_16_0,x[16],y[0]);
and and513(ip_16_1,x[16],y[1]);
and and514(ip_16_2,x[16],y[2]);
and and515(ip_16_3,x[16],y[3]);
and and516(ip_16_4,x[16],y[4]);
and and517(ip_16_5,x[16],y[5]);
and and518(ip_16_6,x[16],y[6]);
and and519(ip_16_7,x[16],y[7]);
and and520(ip_16_8,x[16],y[8]);
and and521(ip_16_9,x[16],y[9]);
and and522(ip_16_10,x[16],y[10]);
and and523(ip_16_11,x[16],y[11]);
and and524(ip_16_12,x[16],y[12]);
and and525(ip_16_13,x[16],y[13]);
and and526(ip_16_14,x[16],y[14]);
and and527(ip_16_15,x[16],y[15]);
and and528(ip_16_16,x[16],y[16]);
and and529(ip_16_17,x[16],y[17]);
and and530(ip_16_18,x[16],y[18]);
and and531(ip_16_19,x[16],y[19]);
and and532(ip_16_20,x[16],y[20]);
and and533(ip_16_21,x[16],y[21]);
and and534(ip_16_22,x[16],y[22]);
and and535(ip_16_23,x[16],y[23]);
and and536(ip_16_24,x[16],y[24]);
and and537(ip_16_25,x[16],y[25]);
and and538(ip_16_26,x[16],y[26]);
and and539(ip_16_27,x[16],y[27]);
and and540(ip_16_28,x[16],y[28]);
and and541(ip_16_29,x[16],y[29]);
and and542(ip_16_30,x[16],y[30]);
and and543(ip_16_31,x[16],y[31]);
and and544(ip_17_0,x[17],y[0]);
and and545(ip_17_1,x[17],y[1]);
and and546(ip_17_2,x[17],y[2]);
and and547(ip_17_3,x[17],y[3]);
and and548(ip_17_4,x[17],y[4]);
and and549(ip_17_5,x[17],y[5]);
and and550(ip_17_6,x[17],y[6]);
and and551(ip_17_7,x[17],y[7]);
and and552(ip_17_8,x[17],y[8]);
and and553(ip_17_9,x[17],y[9]);
and and554(ip_17_10,x[17],y[10]);
and and555(ip_17_11,x[17],y[11]);
and and556(ip_17_12,x[17],y[12]);
and and557(ip_17_13,x[17],y[13]);
and and558(ip_17_14,x[17],y[14]);
and and559(ip_17_15,x[17],y[15]);
and and560(ip_17_16,x[17],y[16]);
and and561(ip_17_17,x[17],y[17]);
and and562(ip_17_18,x[17],y[18]);
and and563(ip_17_19,x[17],y[19]);
and and564(ip_17_20,x[17],y[20]);
and and565(ip_17_21,x[17],y[21]);
and and566(ip_17_22,x[17],y[22]);
and and567(ip_17_23,x[17],y[23]);
and and568(ip_17_24,x[17],y[24]);
and and569(ip_17_25,x[17],y[25]);
and and570(ip_17_26,x[17],y[26]);
and and571(ip_17_27,x[17],y[27]);
and and572(ip_17_28,x[17],y[28]);
and and573(ip_17_29,x[17],y[29]);
and and574(ip_17_30,x[17],y[30]);
and and575(ip_17_31,x[17],y[31]);
and and576(ip_18_0,x[18],y[0]);
and and577(ip_18_1,x[18],y[1]);
and and578(ip_18_2,x[18],y[2]);
and and579(ip_18_3,x[18],y[3]);
and and580(ip_18_4,x[18],y[4]);
and and581(ip_18_5,x[18],y[5]);
and and582(ip_18_6,x[18],y[6]);
and and583(ip_18_7,x[18],y[7]);
and and584(ip_18_8,x[18],y[8]);
and and585(ip_18_9,x[18],y[9]);
and and586(ip_18_10,x[18],y[10]);
and and587(ip_18_11,x[18],y[11]);
and and588(ip_18_12,x[18],y[12]);
and and589(ip_18_13,x[18],y[13]);
and and590(ip_18_14,x[18],y[14]);
and and591(ip_18_15,x[18],y[15]);
and and592(ip_18_16,x[18],y[16]);
and and593(ip_18_17,x[18],y[17]);
and and594(ip_18_18,x[18],y[18]);
and and595(ip_18_19,x[18],y[19]);
and and596(ip_18_20,x[18],y[20]);
and and597(ip_18_21,x[18],y[21]);
and and598(ip_18_22,x[18],y[22]);
and and599(ip_18_23,x[18],y[23]);
and and600(ip_18_24,x[18],y[24]);
and and601(ip_18_25,x[18],y[25]);
and and602(ip_18_26,x[18],y[26]);
and and603(ip_18_27,x[18],y[27]);
and and604(ip_18_28,x[18],y[28]);
and and605(ip_18_29,x[18],y[29]);
and and606(ip_18_30,x[18],y[30]);
and and607(ip_18_31,x[18],y[31]);
and and608(ip_19_0,x[19],y[0]);
and and609(ip_19_1,x[19],y[1]);
and and610(ip_19_2,x[19],y[2]);
and and611(ip_19_3,x[19],y[3]);
and and612(ip_19_4,x[19],y[4]);
and and613(ip_19_5,x[19],y[5]);
and and614(ip_19_6,x[19],y[6]);
and and615(ip_19_7,x[19],y[7]);
and and616(ip_19_8,x[19],y[8]);
and and617(ip_19_9,x[19],y[9]);
and and618(ip_19_10,x[19],y[10]);
and and619(ip_19_11,x[19],y[11]);
and and620(ip_19_12,x[19],y[12]);
and and621(ip_19_13,x[19],y[13]);
and and622(ip_19_14,x[19],y[14]);
and and623(ip_19_15,x[19],y[15]);
and and624(ip_19_16,x[19],y[16]);
and and625(ip_19_17,x[19],y[17]);
and and626(ip_19_18,x[19],y[18]);
and and627(ip_19_19,x[19],y[19]);
and and628(ip_19_20,x[19],y[20]);
and and629(ip_19_21,x[19],y[21]);
and and630(ip_19_22,x[19],y[22]);
and and631(ip_19_23,x[19],y[23]);
and and632(ip_19_24,x[19],y[24]);
and and633(ip_19_25,x[19],y[25]);
and and634(ip_19_26,x[19],y[26]);
and and635(ip_19_27,x[19],y[27]);
and and636(ip_19_28,x[19],y[28]);
and and637(ip_19_29,x[19],y[29]);
and and638(ip_19_30,x[19],y[30]);
and and639(ip_19_31,x[19],y[31]);
and and640(ip_20_0,x[20],y[0]);
and and641(ip_20_1,x[20],y[1]);
and and642(ip_20_2,x[20],y[2]);
and and643(ip_20_3,x[20],y[3]);
and and644(ip_20_4,x[20],y[4]);
and and645(ip_20_5,x[20],y[5]);
and and646(ip_20_6,x[20],y[6]);
and and647(ip_20_7,x[20],y[7]);
and and648(ip_20_8,x[20],y[8]);
and and649(ip_20_9,x[20],y[9]);
and and650(ip_20_10,x[20],y[10]);
and and651(ip_20_11,x[20],y[11]);
and and652(ip_20_12,x[20],y[12]);
and and653(ip_20_13,x[20],y[13]);
and and654(ip_20_14,x[20],y[14]);
and and655(ip_20_15,x[20],y[15]);
and and656(ip_20_16,x[20],y[16]);
and and657(ip_20_17,x[20],y[17]);
and and658(ip_20_18,x[20],y[18]);
and and659(ip_20_19,x[20],y[19]);
and and660(ip_20_20,x[20],y[20]);
and and661(ip_20_21,x[20],y[21]);
and and662(ip_20_22,x[20],y[22]);
and and663(ip_20_23,x[20],y[23]);
and and664(ip_20_24,x[20],y[24]);
and and665(ip_20_25,x[20],y[25]);
and and666(ip_20_26,x[20],y[26]);
and and667(ip_20_27,x[20],y[27]);
and and668(ip_20_28,x[20],y[28]);
and and669(ip_20_29,x[20],y[29]);
and and670(ip_20_30,x[20],y[30]);
and and671(ip_20_31,x[20],y[31]);
and and672(ip_21_0,x[21],y[0]);
and and673(ip_21_1,x[21],y[1]);
and and674(ip_21_2,x[21],y[2]);
and and675(ip_21_3,x[21],y[3]);
and and676(ip_21_4,x[21],y[4]);
and and677(ip_21_5,x[21],y[5]);
and and678(ip_21_6,x[21],y[6]);
and and679(ip_21_7,x[21],y[7]);
and and680(ip_21_8,x[21],y[8]);
and and681(ip_21_9,x[21],y[9]);
and and682(ip_21_10,x[21],y[10]);
and and683(ip_21_11,x[21],y[11]);
and and684(ip_21_12,x[21],y[12]);
and and685(ip_21_13,x[21],y[13]);
and and686(ip_21_14,x[21],y[14]);
and and687(ip_21_15,x[21],y[15]);
and and688(ip_21_16,x[21],y[16]);
and and689(ip_21_17,x[21],y[17]);
and and690(ip_21_18,x[21],y[18]);
and and691(ip_21_19,x[21],y[19]);
and and692(ip_21_20,x[21],y[20]);
and and693(ip_21_21,x[21],y[21]);
and and694(ip_21_22,x[21],y[22]);
and and695(ip_21_23,x[21],y[23]);
and and696(ip_21_24,x[21],y[24]);
and and697(ip_21_25,x[21],y[25]);
and and698(ip_21_26,x[21],y[26]);
and and699(ip_21_27,x[21],y[27]);
and and700(ip_21_28,x[21],y[28]);
and and701(ip_21_29,x[21],y[29]);
and and702(ip_21_30,x[21],y[30]);
and and703(ip_21_31,x[21],y[31]);
and and704(ip_22_0,x[22],y[0]);
and and705(ip_22_1,x[22],y[1]);
and and706(ip_22_2,x[22],y[2]);
and and707(ip_22_3,x[22],y[3]);
and and708(ip_22_4,x[22],y[4]);
and and709(ip_22_5,x[22],y[5]);
and and710(ip_22_6,x[22],y[6]);
and and711(ip_22_7,x[22],y[7]);
and and712(ip_22_8,x[22],y[8]);
and and713(ip_22_9,x[22],y[9]);
and and714(ip_22_10,x[22],y[10]);
and and715(ip_22_11,x[22],y[11]);
and and716(ip_22_12,x[22],y[12]);
and and717(ip_22_13,x[22],y[13]);
and and718(ip_22_14,x[22],y[14]);
and and719(ip_22_15,x[22],y[15]);
and and720(ip_22_16,x[22],y[16]);
and and721(ip_22_17,x[22],y[17]);
and and722(ip_22_18,x[22],y[18]);
and and723(ip_22_19,x[22],y[19]);
and and724(ip_22_20,x[22],y[20]);
and and725(ip_22_21,x[22],y[21]);
and and726(ip_22_22,x[22],y[22]);
and and727(ip_22_23,x[22],y[23]);
and and728(ip_22_24,x[22],y[24]);
and and729(ip_22_25,x[22],y[25]);
and and730(ip_22_26,x[22],y[26]);
and and731(ip_22_27,x[22],y[27]);
and and732(ip_22_28,x[22],y[28]);
and and733(ip_22_29,x[22],y[29]);
and and734(ip_22_30,x[22],y[30]);
and and735(ip_22_31,x[22],y[31]);
and and736(ip_23_0,x[23],y[0]);
and and737(ip_23_1,x[23],y[1]);
and and738(ip_23_2,x[23],y[2]);
and and739(ip_23_3,x[23],y[3]);
and and740(ip_23_4,x[23],y[4]);
and and741(ip_23_5,x[23],y[5]);
and and742(ip_23_6,x[23],y[6]);
and and743(ip_23_7,x[23],y[7]);
and and744(ip_23_8,x[23],y[8]);
and and745(ip_23_9,x[23],y[9]);
and and746(ip_23_10,x[23],y[10]);
and and747(ip_23_11,x[23],y[11]);
and and748(ip_23_12,x[23],y[12]);
and and749(ip_23_13,x[23],y[13]);
and and750(ip_23_14,x[23],y[14]);
and and751(ip_23_15,x[23],y[15]);
and and752(ip_23_16,x[23],y[16]);
and and753(ip_23_17,x[23],y[17]);
and and754(ip_23_18,x[23],y[18]);
and and755(ip_23_19,x[23],y[19]);
and and756(ip_23_20,x[23],y[20]);
and and757(ip_23_21,x[23],y[21]);
and and758(ip_23_22,x[23],y[22]);
and and759(ip_23_23,x[23],y[23]);
and and760(ip_23_24,x[23],y[24]);
and and761(ip_23_25,x[23],y[25]);
and and762(ip_23_26,x[23],y[26]);
and and763(ip_23_27,x[23],y[27]);
and and764(ip_23_28,x[23],y[28]);
and and765(ip_23_29,x[23],y[29]);
and and766(ip_23_30,x[23],y[30]);
and and767(ip_23_31,x[23],y[31]);
and and768(ip_24_0,x[24],y[0]);
and and769(ip_24_1,x[24],y[1]);
and and770(ip_24_2,x[24],y[2]);
and and771(ip_24_3,x[24],y[3]);
and and772(ip_24_4,x[24],y[4]);
and and773(ip_24_5,x[24],y[5]);
and and774(ip_24_6,x[24],y[6]);
and and775(ip_24_7,x[24],y[7]);
and and776(ip_24_8,x[24],y[8]);
and and777(ip_24_9,x[24],y[9]);
and and778(ip_24_10,x[24],y[10]);
and and779(ip_24_11,x[24],y[11]);
and and780(ip_24_12,x[24],y[12]);
and and781(ip_24_13,x[24],y[13]);
and and782(ip_24_14,x[24],y[14]);
and and783(ip_24_15,x[24],y[15]);
and and784(ip_24_16,x[24],y[16]);
and and785(ip_24_17,x[24],y[17]);
and and786(ip_24_18,x[24],y[18]);
and and787(ip_24_19,x[24],y[19]);
and and788(ip_24_20,x[24],y[20]);
and and789(ip_24_21,x[24],y[21]);
and and790(ip_24_22,x[24],y[22]);
and and791(ip_24_23,x[24],y[23]);
and and792(ip_24_24,x[24],y[24]);
and and793(ip_24_25,x[24],y[25]);
and and794(ip_24_26,x[24],y[26]);
and and795(ip_24_27,x[24],y[27]);
and and796(ip_24_28,x[24],y[28]);
and and797(ip_24_29,x[24],y[29]);
and and798(ip_24_30,x[24],y[30]);
and and799(ip_24_31,x[24],y[31]);
and and800(ip_25_0,x[25],y[0]);
and and801(ip_25_1,x[25],y[1]);
and and802(ip_25_2,x[25],y[2]);
and and803(ip_25_3,x[25],y[3]);
and and804(ip_25_4,x[25],y[4]);
and and805(ip_25_5,x[25],y[5]);
and and806(ip_25_6,x[25],y[6]);
and and807(ip_25_7,x[25],y[7]);
and and808(ip_25_8,x[25],y[8]);
and and809(ip_25_9,x[25],y[9]);
and and810(ip_25_10,x[25],y[10]);
and and811(ip_25_11,x[25],y[11]);
and and812(ip_25_12,x[25],y[12]);
and and813(ip_25_13,x[25],y[13]);
and and814(ip_25_14,x[25],y[14]);
and and815(ip_25_15,x[25],y[15]);
and and816(ip_25_16,x[25],y[16]);
and and817(ip_25_17,x[25],y[17]);
and and818(ip_25_18,x[25],y[18]);
and and819(ip_25_19,x[25],y[19]);
and and820(ip_25_20,x[25],y[20]);
and and821(ip_25_21,x[25],y[21]);
and and822(ip_25_22,x[25],y[22]);
and and823(ip_25_23,x[25],y[23]);
and and824(ip_25_24,x[25],y[24]);
and and825(ip_25_25,x[25],y[25]);
and and826(ip_25_26,x[25],y[26]);
and and827(ip_25_27,x[25],y[27]);
and and828(ip_25_28,x[25],y[28]);
and and829(ip_25_29,x[25],y[29]);
and and830(ip_25_30,x[25],y[30]);
and and831(ip_25_31,x[25],y[31]);
and and832(ip_26_0,x[26],y[0]);
and and833(ip_26_1,x[26],y[1]);
and and834(ip_26_2,x[26],y[2]);
and and835(ip_26_3,x[26],y[3]);
and and836(ip_26_4,x[26],y[4]);
and and837(ip_26_5,x[26],y[5]);
and and838(ip_26_6,x[26],y[6]);
and and839(ip_26_7,x[26],y[7]);
and and840(ip_26_8,x[26],y[8]);
and and841(ip_26_9,x[26],y[9]);
and and842(ip_26_10,x[26],y[10]);
and and843(ip_26_11,x[26],y[11]);
and and844(ip_26_12,x[26],y[12]);
and and845(ip_26_13,x[26],y[13]);
and and846(ip_26_14,x[26],y[14]);
and and847(ip_26_15,x[26],y[15]);
and and848(ip_26_16,x[26],y[16]);
and and849(ip_26_17,x[26],y[17]);
and and850(ip_26_18,x[26],y[18]);
and and851(ip_26_19,x[26],y[19]);
and and852(ip_26_20,x[26],y[20]);
and and853(ip_26_21,x[26],y[21]);
and and854(ip_26_22,x[26],y[22]);
and and855(ip_26_23,x[26],y[23]);
and and856(ip_26_24,x[26],y[24]);
and and857(ip_26_25,x[26],y[25]);
and and858(ip_26_26,x[26],y[26]);
and and859(ip_26_27,x[26],y[27]);
and and860(ip_26_28,x[26],y[28]);
and and861(ip_26_29,x[26],y[29]);
and and862(ip_26_30,x[26],y[30]);
and and863(ip_26_31,x[26],y[31]);
and and864(ip_27_0,x[27],y[0]);
and and865(ip_27_1,x[27],y[1]);
and and866(ip_27_2,x[27],y[2]);
and and867(ip_27_3,x[27],y[3]);
and and868(ip_27_4,x[27],y[4]);
and and869(ip_27_5,x[27],y[5]);
and and870(ip_27_6,x[27],y[6]);
and and871(ip_27_7,x[27],y[7]);
and and872(ip_27_8,x[27],y[8]);
and and873(ip_27_9,x[27],y[9]);
and and874(ip_27_10,x[27],y[10]);
and and875(ip_27_11,x[27],y[11]);
and and876(ip_27_12,x[27],y[12]);
and and877(ip_27_13,x[27],y[13]);
and and878(ip_27_14,x[27],y[14]);
and and879(ip_27_15,x[27],y[15]);
and and880(ip_27_16,x[27],y[16]);
and and881(ip_27_17,x[27],y[17]);
and and882(ip_27_18,x[27],y[18]);
and and883(ip_27_19,x[27],y[19]);
and and884(ip_27_20,x[27],y[20]);
and and885(ip_27_21,x[27],y[21]);
and and886(ip_27_22,x[27],y[22]);
and and887(ip_27_23,x[27],y[23]);
and and888(ip_27_24,x[27],y[24]);
and and889(ip_27_25,x[27],y[25]);
and and890(ip_27_26,x[27],y[26]);
and and891(ip_27_27,x[27],y[27]);
and and892(ip_27_28,x[27],y[28]);
and and893(ip_27_29,x[27],y[29]);
and and894(ip_27_30,x[27],y[30]);
and and895(ip_27_31,x[27],y[31]);
and and896(ip_28_0,x[28],y[0]);
and and897(ip_28_1,x[28],y[1]);
and and898(ip_28_2,x[28],y[2]);
and and899(ip_28_3,x[28],y[3]);
and and900(ip_28_4,x[28],y[4]);
and and901(ip_28_5,x[28],y[5]);
and and902(ip_28_6,x[28],y[6]);
and and903(ip_28_7,x[28],y[7]);
and and904(ip_28_8,x[28],y[8]);
and and905(ip_28_9,x[28],y[9]);
and and906(ip_28_10,x[28],y[10]);
and and907(ip_28_11,x[28],y[11]);
and and908(ip_28_12,x[28],y[12]);
and and909(ip_28_13,x[28],y[13]);
and and910(ip_28_14,x[28],y[14]);
and and911(ip_28_15,x[28],y[15]);
and and912(ip_28_16,x[28],y[16]);
and and913(ip_28_17,x[28],y[17]);
and and914(ip_28_18,x[28],y[18]);
and and915(ip_28_19,x[28],y[19]);
and and916(ip_28_20,x[28],y[20]);
and and917(ip_28_21,x[28],y[21]);
and and918(ip_28_22,x[28],y[22]);
and and919(ip_28_23,x[28],y[23]);
and and920(ip_28_24,x[28],y[24]);
and and921(ip_28_25,x[28],y[25]);
and and922(ip_28_26,x[28],y[26]);
and and923(ip_28_27,x[28],y[27]);
and and924(ip_28_28,x[28],y[28]);
and and925(ip_28_29,x[28],y[29]);
and and926(ip_28_30,x[28],y[30]);
and and927(ip_28_31,x[28],y[31]);
and and928(ip_29_0,x[29],y[0]);
and and929(ip_29_1,x[29],y[1]);
and and930(ip_29_2,x[29],y[2]);
and and931(ip_29_3,x[29],y[3]);
and and932(ip_29_4,x[29],y[4]);
and and933(ip_29_5,x[29],y[5]);
and and934(ip_29_6,x[29],y[6]);
and and935(ip_29_7,x[29],y[7]);
and and936(ip_29_8,x[29],y[8]);
and and937(ip_29_9,x[29],y[9]);
and and938(ip_29_10,x[29],y[10]);
and and939(ip_29_11,x[29],y[11]);
and and940(ip_29_12,x[29],y[12]);
and and941(ip_29_13,x[29],y[13]);
and and942(ip_29_14,x[29],y[14]);
and and943(ip_29_15,x[29],y[15]);
and and944(ip_29_16,x[29],y[16]);
and and945(ip_29_17,x[29],y[17]);
and and946(ip_29_18,x[29],y[18]);
and and947(ip_29_19,x[29],y[19]);
and and948(ip_29_20,x[29],y[20]);
and and949(ip_29_21,x[29],y[21]);
and and950(ip_29_22,x[29],y[22]);
and and951(ip_29_23,x[29],y[23]);
and and952(ip_29_24,x[29],y[24]);
and and953(ip_29_25,x[29],y[25]);
and and954(ip_29_26,x[29],y[26]);
and and955(ip_29_27,x[29],y[27]);
and and956(ip_29_28,x[29],y[28]);
and and957(ip_29_29,x[29],y[29]);
and and958(ip_29_30,x[29],y[30]);
and and959(ip_29_31,x[29],y[31]);
and and960(ip_30_0,x[30],y[0]);
and and961(ip_30_1,x[30],y[1]);
and and962(ip_30_2,x[30],y[2]);
and and963(ip_30_3,x[30],y[3]);
and and964(ip_30_4,x[30],y[4]);
and and965(ip_30_5,x[30],y[5]);
and and966(ip_30_6,x[30],y[6]);
and and967(ip_30_7,x[30],y[7]);
and and968(ip_30_8,x[30],y[8]);
and and969(ip_30_9,x[30],y[9]);
and and970(ip_30_10,x[30],y[10]);
and and971(ip_30_11,x[30],y[11]);
and and972(ip_30_12,x[30],y[12]);
and and973(ip_30_13,x[30],y[13]);
and and974(ip_30_14,x[30],y[14]);
and and975(ip_30_15,x[30],y[15]);
and and976(ip_30_16,x[30],y[16]);
and and977(ip_30_17,x[30],y[17]);
and and978(ip_30_18,x[30],y[18]);
and and979(ip_30_19,x[30],y[19]);
and and980(ip_30_20,x[30],y[20]);
and and981(ip_30_21,x[30],y[21]);
and and982(ip_30_22,x[30],y[22]);
and and983(ip_30_23,x[30],y[23]);
and and984(ip_30_24,x[30],y[24]);
and and985(ip_30_25,x[30],y[25]);
and and986(ip_30_26,x[30],y[26]);
and and987(ip_30_27,x[30],y[27]);
and and988(ip_30_28,x[30],y[28]);
and and989(ip_30_29,x[30],y[29]);
and and990(ip_30_30,x[30],y[30]);
and and991(ip_30_31,x[30],y[31]);
and and992(ip_31_0,x[31],y[0]);
and and993(ip_31_1,x[31],y[1]);
and and994(ip_31_2,x[31],y[2]);
and and995(ip_31_3,x[31],y[3]);
and and996(ip_31_4,x[31],y[4]);
and and997(ip_31_5,x[31],y[5]);
and and998(ip_31_6,x[31],y[6]);
and and999(ip_31_7,x[31],y[7]);
and and1000(ip_31_8,x[31],y[8]);
and and1001(ip_31_9,x[31],y[9]);
and and1002(ip_31_10,x[31],y[10]);
and and1003(ip_31_11,x[31],y[11]);
and and1004(ip_31_12,x[31],y[12]);
and and1005(ip_31_13,x[31],y[13]);
and and1006(ip_31_14,x[31],y[14]);
and and1007(ip_31_15,x[31],y[15]);
and and1008(ip_31_16,x[31],y[16]);
and and1009(ip_31_17,x[31],y[17]);
and and1010(ip_31_18,x[31],y[18]);
and and1011(ip_31_19,x[31],y[19]);
and and1012(ip_31_20,x[31],y[20]);
and and1013(ip_31_21,x[31],y[21]);
and and1014(ip_31_22,x[31],y[22]);
and and1015(ip_31_23,x[31],y[23]);
and and1016(ip_31_24,x[31],y[24]);
and and1017(ip_31_25,x[31],y[25]);
and and1018(ip_31_26,x[31],y[26]);
and and1019(ip_31_27,x[31],y[27]);
and and1020(ip_31_28,x[31],y[28]);
and and1021(ip_31_29,x[31],y[29]);
and and1022(ip_31_30,x[31],y[30]);
and and1023(ip_31_31,x[31],y[31]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
HA ha0(ip_3_0,p3,p4,p5);
HA ha1(ip_0_4,ip_1_3,p6,p7);
FA fa2(ip_2_2,ip_3_1,ip_4_0,p8,p9);
FA fa3(p7,p9,p2,p10,p11);
FA fa4(ip_0_5,ip_1_4,ip_2_3,p12,p13);
FA fa5(ip_3_2,ip_4_1,ip_5_0,p14,p15);
FA fa6(p6,p13,p15,p16,p17);
FA fa7(p8,p17,p10,p18,p19);
HA ha2(ip_0_6,ip_1_5,p20,p21);
HA ha3(ip_2_4,ip_3_3,p22,p23);
HA ha4(ip_4_2,ip_5_1,p24,p25);
HA ha5(ip_6_0,p21,p26,p27);
FA fa8(p23,p25,p27,p28,p29);
FA fa9(p12,p14,p29,p30,p31);
HA ha6(p16,p31,p32,p33);
HA ha7(ip_0_7,ip_1_6,p34,p35);
FA fa10(ip_2_5,ip_3_4,ip_4_3,p36,p37);
FA fa11(ip_5_2,ip_6_1,ip_7_0,p38,p39);
FA fa12(p20,p22,p24,p40,p41);
HA ha8(p35,p26,p42,p43);
HA ha9(p37,p39,p44,p45);
HA ha10(p41,p43,p46,p47);
FA fa13(p45,p28,p47,p48,p49);
HA ha11(p30,p32,p50,p51);
FA fa14(ip_0_8,ip_1_7,ip_2_6,p52,p53);
HA ha12(ip_3_5,ip_4_4,p54,p55);
FA fa15(ip_5_3,ip_6_2,ip_7_1,p56,p57);
FA fa16(ip_8_0,p34,p55,p58,p59);
HA ha13(p53,p57,p60,p61);
FA fa17(p36,p38,p42,p62,p63);
FA fa18(p44,p59,p61,p64,p65);
HA ha14(p40,p46,p66,p67);
HA ha15(p63,p65,p68,p69);
FA fa19(p67,p69,p48,p70,p71);
FA fa20(ip_0_9,ip_1_8,ip_2_7,p72,p73);
HA ha16(ip_3_6,ip_4_5,p74,p75);
HA ha17(ip_5_4,ip_6_3,p76,p77);
HA ha18(ip_7_2,ip_8_1,p78,p79);
HA ha19(ip_9_0,p54,p80,p81);
FA fa21(p75,p77,p79,p82,p83);
FA fa22(p73,p81,p52,p84,p85);
FA fa23(p56,p60,p83,p86,p87);
FA fa24(p58,p85,p66,p88,p89);
HA ha20(p87,p62,p90,p91);
FA fa25(p64,p68,p89,p92,p93);
FA fa26(p91,p93,p70,p94,p95);
FA fa27(ip_0_10,ip_1_9,ip_2_8,p96,p97);
HA ha21(ip_3_7,ip_4_6,p98,p99);
FA fa28(ip_5_5,ip_6_4,ip_7_3,p100,p101);
HA ha22(ip_8_2,ip_9_1,p102,p103);
FA fa29(ip_10_0,p103,p74,p104,p105);
HA ha23(p76,p78,p106,p107);
HA ha24(p99,p101,p108,p109);
FA fa30(p107,p80,p97,p110,p111);
FA fa31(p105,p109,p72,p112,p113);
FA fa32(p111,p82,p113,p114,p115);
FA fa33(p84,p115,p86,p116,p117);
FA fa34(p88,p90,p117,p118,p119);
HA ha25(p119,p92,p120,p121);
FA fa35(ip_0_11,ip_1_10,ip_2_9,p122,p123);
FA fa36(ip_3_8,ip_4_7,ip_5_6,p124,p125);
FA fa37(ip_6_5,ip_7_4,ip_8_3,p126,p127);
HA ha26(ip_9_2,ip_10_1,p128,p129);
HA ha27(ip_11_0,p102,p130,p131);
HA ha28(p129,p98,p132,p133);
HA ha29(p106,p123,p134,p135);
FA fa38(p125,p127,p131,p136,p137);
FA fa39(p133,p100,p108,p138,p139);
FA fa40(p135,p96,p104,p140,p141);
HA ha30(p137,p110,p142,p143);
FA fa41(p139,p141,p112,p144,p145);
FA fa42(p143,p114,p145,p146,p147);
FA fa43(p116,p147,p118,p148,p149);
HA ha31(ip_0_12,ip_1_11,p150,p151);
FA fa44(ip_2_10,ip_3_9,ip_4_8,p152,p153);
FA fa45(ip_5_7,ip_6_6,ip_7_5,p154,p155);
FA fa46(ip_8_4,ip_9_3,ip_10_2,p156,p157);
HA ha32(ip_11_1,ip_12_0,p158,p159);
HA ha33(p128,p151,p160,p161);
HA ha34(p159,p130,p162,p163);
FA fa47(p132,p153,p155,p164,p165);
HA ha35(p157,p161,p166,p167);
FA fa48(p122,p124,p126,p168,p169);
FA fa49(p134,p163,p167,p170,p171);
FA fa50(p165,p136,p169,p172,p173);
FA fa51(p171,p138,p140,p174,p175);
HA ha36(p142,p173,p176,p177);
FA fa52(p144,p175,p177,p178,p179);
HA ha37(p146,p179,p180,p181);
HA ha38(ip_0_13,ip_1_12,p182,p183);
HA ha39(ip_2_11,ip_3_10,p184,p185);
HA ha40(ip_4_9,ip_5_8,p186,p187);
FA fa53(ip_6_7,ip_7_6,ip_8_5,p188,p189);
HA ha41(ip_9_4,ip_10_3,p190,p191);
HA ha42(ip_11_2,ip_12_1,p192,p193);
FA fa54(ip_13_0,p150,p158,p194,p195);
FA fa55(p183,p185,p187,p196,p197);
FA fa56(p191,p193,p160,p198,p199);
HA ha43(p189,p152,p200,p201);
HA ha44(p154,p156,p202,p203);
FA fa57(p162,p166,p195,p204,p205);
HA ha45(p197,p199,p206,p207);
FA fa58(p201,p203,p207,p208,p209);
FA fa59(p164,p205,p168,p210,p211);
HA ha46(p170,p209,p212,p213);
FA fa60(p211,p213,p172,p214,p215);
HA ha47(p176,p174,p216,p217);
HA ha48(p215,p217,p218,p219);
HA ha49(p178,p180,p220,p221);
HA ha50(ip_0_14,ip_1_13,p222,p223);
FA fa61(ip_2_12,ip_3_11,ip_4_10,p224,p225);
FA fa62(ip_5_9,ip_6_8,ip_7_7,p226,p227);
FA fa63(ip_8_6,ip_9_5,ip_10_4,p228,p229);
HA ha51(ip_11_3,ip_12_2,p230,p231);
HA ha52(ip_13_1,ip_14_0,p232,p233);
HA ha53(p182,p184,p234,p235);
HA ha54(p186,p190,p236,p237);
HA ha55(p192,p223,p238,p239);
FA fa64(p231,p233,p225,p240,p241);
FA fa65(p227,p229,p235,p242,p243);
HA ha56(p237,p239,p244,p245);
HA ha57(p188,p241,p246,p247);
FA fa66(p245,p194,p196,p248,p249);
FA fa67(p198,p200,p202,p250,p251);
FA fa68(p206,p243,p247,p252,p253);
HA ha58(p204,p249,p254,p255);
HA ha59(p251,p253,p256,p257);
HA ha60(p208,p212,p258,p259);
FA fa69(p255,p257,p210,p260,p261);
FA fa70(p259,p261,p214,p262,p263);
HA ha61(p216,p218,p264,p265);
HA ha62(p263,p220,p266,p267);
FA fa71(ip_0_15,ip_1_14,ip_2_13,p268,p269);
HA ha63(ip_3_12,ip_4_11,p270,p271);
FA fa72(ip_5_10,ip_6_9,ip_7_8,p272,p273);
FA fa73(ip_8_7,ip_9_6,ip_10_5,p274,p275);
HA ha64(ip_11_4,ip_12_3,p276,p277);
FA fa74(ip_13_2,ip_14_1,ip_15_0,p278,p279);
FA fa75(p222,p230,p232,p280,p281);
HA ha65(p271,p277,p282,p283);
HA ha66(p234,p236,p284,p285);
FA fa76(p238,p269,p273,p286,p287);
HA ha67(p275,p279,p288,p289);
HA ha68(p283,p224,p290,p291);
FA fa77(p226,p228,p244,p292,p293);
FA fa78(p281,p285,p289,p294,p295);
HA ha69(p240,p246,p296,p297);
HA ha70(p287,p291,p298,p299);
FA fa79(p242,p293,p295,p300,p301);
HA ha71(p297,p299,p302,p303);
FA fa80(p303,p248,p250,p304,p305);
FA fa81(p252,p254,p256,p306,p307);
HA ha72(p301,p258,p308,p309);
HA ha73(p305,p307,p310,p311);
HA ha74(p309,p260,p312,p313);
FA fa82(p311,p313,p262,p314,p315);
HA ha75(p264,p266,p316,p317);
FA fa83(ip_0_16,ip_1_15,ip_2_14,p318,p319);
HA ha76(ip_3_13,ip_4_12,p320,p321);
FA fa84(ip_5_11,ip_6_10,ip_7_9,p322,p323);
FA fa85(ip_8_8,ip_9_7,ip_10_6,p324,p325);
HA ha77(ip_11_5,ip_12_4,p326,p327);
FA fa86(ip_13_3,ip_14_2,ip_15_1,p328,p329);
HA ha78(ip_16_0,p270,p330,p331);
HA ha79(p276,p321,p332,p333);
HA ha80(p327,p282,p334,p335);
FA fa87(p319,p323,p325,p336,p337);
HA ha81(p329,p331,p338,p339);
FA fa88(p333,p268,p272,p340,p341);
FA fa89(p274,p278,p284,p342,p343);
HA ha82(p288,p335,p344,p345);
HA ha83(p339,p280,p346,p347);
HA ha84(p290,p337,p348,p349);
FA fa90(p345,p286,p296,p350,p351);
HA ha85(p298,p341,p352,p353);
HA ha86(p343,p347,p354,p355);
HA ha87(p349,p292,p356,p357);
FA fa91(p294,p302,p353,p358,p359);
HA ha88(p355,p351,p360,p361);
FA fa92(p357,p300,p359,p362,p363);
FA fa93(p361,p308,p304,p364,p365);
FA fa94(p306,p310,p363,p366,p367);
HA ha89(p312,p365,p368,p369);
HA ha90(p367,p369,p370,p371);
FA fa95(p371,p314,p316,p372,p373);
FA fa96(ip_0_17,ip_1_16,ip_2_15,p374,p375);
HA ha91(ip_3_14,ip_4_13,p376,p377);
HA ha92(ip_5_12,ip_6_11,p378,p379);
FA fa97(ip_7_10,ip_8_9,ip_9_8,p380,p381);
HA ha93(ip_10_7,ip_11_6,p382,p383);
HA ha94(ip_12_5,ip_13_4,p384,p385);
FA fa98(ip_14_3,ip_15_2,ip_16_1,p386,p387);
HA ha95(ip_17_0,p320,p388,p389);
FA fa99(p326,p377,p379,p390,p391);
FA fa100(p383,p385,p330,p392,p393);
FA fa101(p332,p375,p381,p394,p395);
FA fa102(p387,p389,p318,p396,p397);
FA fa103(p322,p324,p328,p398,p399);
FA fa104(p334,p338,p391,p400,p401);
FA fa105(p393,p344,p395,p402,p403);
HA ha96(p397,p336,p404,p405);
HA ha97(p346,p348,p406,p407);
HA ha98(p399,p401,p408,p409);
FA fa106(p340,p342,p352,p410,p411);
FA fa107(p354,p403,p405,p412,p413);
FA fa108(p407,p409,p356,p414,p415);
HA ha99(p350,p360,p416,p417);
FA fa109(p411,p413,p415,p418,p419);
FA fa110(p358,p417,p419,p420,p421);
HA ha100(p362,p421,p422,p423);
FA fa111(p364,p368,p423,p424,p425);
HA ha101(p366,p370,p426,p427);
FA fa112(p425,p427,p372,p428,p429);
HA ha102(ip_0_18,ip_1_17,p430,p431);
HA ha103(ip_2_16,ip_3_15,p432,p433);
HA ha104(ip_4_14,ip_5_13,p434,p435);
HA ha105(ip_6_12,ip_7_11,p436,p437);
FA fa113(ip_8_10,ip_9_9,ip_10_8,p438,p439);
HA ha106(ip_11_7,ip_12_6,p440,p441);
HA ha107(ip_13_5,ip_14_4,p442,p443);
FA fa114(ip_15_3,ip_16_2,ip_17_1,p444,p445);
FA fa115(ip_18_0,p376,p378,p446,p447);
HA ha108(p382,p384,p448,p449);
HA ha109(p431,p433,p450,p451);
FA fa116(p435,p437,p441,p452,p453);
FA fa117(p443,p388,p439,p454,p455);
HA ha110(p445,p449,p456,p457);
HA ha111(p451,p374,p458,p459);
FA fa118(p380,p386,p447,p460,p461);
FA fa119(p453,p457,p390,p462,p463);
FA fa120(p392,p455,p459,p464,p465);
FA fa121(p394,p396,p461,p466,p467);
FA fa122(p463,p398,p400,p468,p469);
HA ha112(p404,p406,p470,p471);
HA ha113(p408,p465,p472,p473);
HA ha114(p402,p467,p474,p475);
FA fa123(p471,p473,p469,p476,p477);
FA fa124(p475,p410,p412,p478,p479);
HA ha115(p414,p416,p480,p481);
HA ha116(p477,p481,p482,p483);
FA fa125(p418,p479,p483,p484,p485);
FA fa126(p420,p422,p485,p486,p487);
HA ha117(p426,p487,p488,p489);
FA fa127(p424,p489,p428,p490,p491);
FA fa128(ip_0_19,ip_1_18,ip_2_17,p492,p493);
FA fa129(ip_3_16,ip_4_15,ip_5_14,p494,p495);
HA ha118(ip_6_13,ip_7_12,p496,p497);
FA fa130(ip_8_11,ip_9_10,ip_10_9,p498,p499);
FA fa131(ip_11_8,ip_12_7,ip_13_6,p500,p501);
HA ha119(ip_14_5,ip_15_4,p502,p503);
FA fa132(ip_16_3,ip_17_2,ip_18_1,p504,p505);
FA fa133(ip_19_0,p430,p432,p506,p507);
FA fa134(p434,p436,p440,p508,p509);
HA ha120(p442,p497,p510,p511);
FA fa135(p503,p448,p450,p512,p513);
HA ha121(p493,p495,p514,p515);
FA fa136(p499,p501,p505,p516,p517);
FA fa137(p511,p438,p444,p518,p519);
HA ha122(p456,p507,p520,p521);
FA fa138(p509,p515,p446,p522,p523);
HA ha123(p452,p458,p524,p525);
HA ha124(p513,p517,p526,p527);
HA ha125(p521,p454,p528,p529);
HA ha126(p519,p523,p530,p531);
FA fa139(p525,p527,p460,p532,p533);
FA fa140(p462,p529,p531,p534,p535);
FA fa141(p464,p470,p472,p536,p537);
HA ha127(p533,p466,p538,p539);
FA fa142(p474,p535,p468,p540,p541);
FA fa143(p537,p539,p476,p542,p543);
FA fa144(p480,p541,p482,p544,p545);
HA ha128(p543,p478,p546,p547);
FA fa145(p545,p547,p484,p548,p549);
FA fa146(p486,p488,p549,p550,p551);
HA ha129(ip_0_20,ip_1_19,p552,p553);
FA fa147(ip_2_18,ip_3_17,ip_4_16,p554,p555);
HA ha130(ip_5_15,ip_6_14,p556,p557);
FA fa148(ip_7_13,ip_8_12,ip_9_11,p558,p559);
FA fa149(ip_10_10,ip_11_9,ip_12_8,p560,p561);
HA ha131(ip_13_7,ip_14_6,p562,p563);
FA fa150(ip_15_5,ip_16_4,ip_17_3,p564,p565);
FA fa151(ip_18_2,ip_19_1,ip_20_0,p566,p567);
HA ha132(p496,p502,p568,p569);
HA ha133(p553,p557,p570,p571);
FA fa152(p563,p510,p555,p572,p573);
FA fa153(p559,p561,p565,p574,p575);
HA ha134(p567,p569,p576,p577);
FA fa154(p571,p492,p494,p578,p579);
HA ha135(p498,p500,p580,p581);
HA ha136(p504,p514,p582,p583);
HA ha137(p577,p506,p584,p585);
HA ha138(p508,p520,p586,p587);
FA fa155(p573,p575,p581,p588,p589);
HA ha139(p583,p512,p590,p591);
FA fa156(p516,p524,p526,p592,p593);
FA fa157(p579,p585,p587,p594,p595);
HA ha140(p518,p522,p596,p597);
HA ha141(p528,p530,p598,p599);
HA ha142(p589,p591,p600,p601);
FA fa158(p593,p595,p597,p602,p603);
HA ha143(p599,p601,p604,p605);
FA fa159(p532,p605,p534,p606,p607);
FA fa160(p538,p603,p536,p608,p609);
HA ha144(p607,p540,p610,p611);
HA ha145(p609,p542,p612,p613);
HA ha146(p611,p544,p614,p615);
FA fa161(p546,p613,p615,p616,p617);
HA ha147(p617,p548,p618,p619);
FA fa162(ip_0_21,ip_1_20,ip_2_19,p620,p621);
HA ha148(ip_3_18,ip_4_17,p622,p623);
FA fa163(ip_5_16,ip_6_15,ip_7_14,p624,p625);
HA ha149(ip_8_13,ip_9_12,p626,p627);
HA ha150(ip_10_11,ip_11_10,p628,p629);
FA fa164(ip_12_9,ip_13_8,ip_14_7,p630,p631);
HA ha151(ip_15_6,ip_16_5,p632,p633);
FA fa165(ip_17_4,ip_18_3,ip_19_2,p634,p635);
FA fa166(ip_20_1,ip_21_0,p552,p636,p637);
HA ha152(p556,p562,p638,p639);
FA fa167(p623,p627,p629,p640,p641);
FA fa168(p633,p568,p570,p642,p643);
FA fa169(p621,p625,p631,p644,p645);
FA fa170(p635,p637,p639,p646,p647);
HA ha153(p554,p558,p648,p649);
HA ha154(p560,p564,p650,p651);
FA fa171(p566,p576,p641,p652,p653);
FA fa172(p580,p582,p643,p654,p655);
FA fa173(p645,p647,p649,p656,p657);
HA ha155(p651,p572,p658,p659);
HA ha156(p574,p584,p660,p661);
FA fa174(p586,p653,p578,p662,p663);
FA fa175(p590,p655,p657,p664,p665);
FA fa176(p659,p661,p588,p666,p667);
FA fa177(p596,p598,p600,p668,p669);
FA fa178(p663,p592,p594,p670,p671);
HA ha157(p604,p665,p672,p673);
FA fa179(p667,p669,p673,p674,p675);
FA fa180(p602,p671,p606,p676,p677);
HA ha158(p675,p608,p678,p679);
HA ha159(p610,p677,p680,p681);
HA ha160(p612,p679,p682,p683);
FA fa181(p681,p614,p683,p684,p685);
HA ha161(p616,p685,p686,p687);
HA ha162(ip_0_22,ip_1_21,p688,p689);
FA fa182(ip_2_20,ip_3_19,ip_4_18,p690,p691);
HA ha163(ip_5_17,ip_6_16,p692,p693);
FA fa183(ip_7_15,ip_8_14,ip_9_13,p694,p695);
FA fa184(ip_10_12,ip_11_11,ip_12_10,p696,p697);
FA fa185(ip_13_9,ip_14_8,ip_15_7,p698,p699);
HA ha164(ip_16_6,ip_17_5,p700,p701);
FA fa186(ip_18_4,ip_19_3,ip_20_2,p702,p703);
FA fa187(ip_21_1,ip_22_0,p622,p704,p705);
HA ha165(p626,p628,p706,p707);
FA fa188(p632,p689,p693,p708,p709);
FA fa189(p701,p638,p691,p710,p711);
FA fa190(p695,p697,p699,p712,p713);
FA fa191(p703,p705,p707,p714,p715);
HA ha166(p620,p624,p716,p717);
HA ha167(p630,p634,p718,p719);
HA ha168(p636,p709,p720,p721);
HA ha169(p640,p648,p722,p723);
HA ha170(p650,p711,p724,p725);
HA ha171(p713,p715,p726,p727);
FA fa192(p717,p719,p721,p728,p729);
HA ha172(p642,p644,p730,p731);
HA ha173(p646,p723,p732,p733);
FA fa193(p725,p727,p652,p734,p735);
FA fa194(p658,p660,p729,p736,p737);
HA ha174(p731,p733,p738,p739);
HA ha175(p654,p656,p740,p741);
HA ha176(p735,p739,p742,p743);
HA ha177(p662,p737,p744,p745);
HA ha178(p741,p743,p746,p747);
HA ha179(p664,p666,p748,p749);
FA fa195(p672,p745,p747,p750,p751);
HA ha180(p668,p749,p752,p753);
FA fa196(p670,p751,p753,p754,p755);
HA ha181(p674,p676,p756,p757);
FA fa197(p678,p680,p755,p758,p759);
FA fa198(p682,p757,p759,p760,p761);
FA fa199(p761,p684,p686,p762,p763);
HA ha182(ip_0_23,ip_1_22,p764,p765);
FA fa200(ip_2_21,ip_3_20,ip_4_19,p766,p767);
HA ha183(ip_5_18,ip_6_17,p768,p769);
HA ha184(ip_7_16,ip_8_15,p770,p771);
FA fa201(ip_9_14,ip_10_13,ip_11_12,p772,p773);
HA ha185(ip_12_11,ip_13_10,p774,p775);
HA ha186(ip_14_9,ip_15_8,p776,p777);
HA ha187(ip_16_7,ip_17_6,p778,p779);
FA fa202(ip_18_5,ip_19_4,ip_20_3,p780,p781);
HA ha188(ip_21_2,ip_22_1,p782,p783);
HA ha189(ip_23_0,p688,p784,p785);
FA fa203(p692,p700,p765,p786,p787);
FA fa204(p769,p771,p775,p788,p789);
HA ha190(p777,p779,p790,p791);
HA ha191(p783,p706,p792,p793);
HA ha192(p767,p773,p794,p795);
FA fa205(p781,p785,p791,p796,p797);
HA ha193(p690,p694,p798,p799);
HA ha194(p696,p698,p800,p801);
HA ha195(p702,p704,p802,p803);
HA ha196(p787,p789,p804,p805);
FA fa206(p793,p795,p708,p806,p807);
FA fa207(p716,p718,p720,p808,p809);
HA ha197(p797,p799,p810,p811);
FA fa208(p801,p803,p805,p812,p813);
FA fa209(p710,p712,p714,p814,p815);
HA ha198(p722,p724,p816,p817);
HA ha199(p726,p807,p818,p819);
HA ha200(p811,p730,p820,p821);
HA ha201(p732,p809,p822,p823);
FA fa210(p813,p817,p819,p824,p825);
FA fa211(p728,p738,p815,p826,p827);
FA fa212(p821,p823,p734,p828,p829);
HA ha202(p740,p742,p830,p831);
FA fa213(p825,p736,p744,p832,p833);
HA ha203(p746,p827,p834,p835);
HA ha204(p829,p831,p836,p837);
FA fa214(p748,p835,p837,p838,p839);
HA ha205(p752,p833,p840,p841);
HA ha206(p750,p839,p842,p843);
FA fa215(p841,p843,p754,p844,p845);
FA fa216(p756,p845,p758,p846,p847);
HA ha207(p760,p847,p848,p849);
FA fa217(ip_0_24,ip_1_23,ip_2_22,p850,p851);
FA fa218(ip_3_21,ip_4_20,ip_5_19,p852,p853);
FA fa219(ip_6_18,ip_7_17,ip_8_16,p854,p855);
FA fa220(ip_9_15,ip_10_14,ip_11_13,p856,p857);
HA ha208(ip_12_12,ip_13_11,p858,p859);
HA ha209(ip_14_10,ip_15_9,p860,p861);
FA fa221(ip_16_8,ip_17_7,ip_18_6,p862,p863);
FA fa222(ip_19_5,ip_20_4,ip_21_3,p864,p865);
HA ha210(ip_22_2,ip_23_1,p866,p867);
HA ha211(ip_24_0,p764,p868,p869);
HA ha212(p768,p770,p870,p871);
FA fa223(p774,p776,p778,p872,p873);
HA ha213(p782,p859,p874,p875);
FA fa224(p861,p867,p784,p876,p877);
FA fa225(p790,p851,p853,p878,p879);
HA ha214(p855,p857,p880,p881);
HA ha215(p863,p865,p882,p883);
FA fa226(p869,p871,p875,p884,p885);
FA fa227(p766,p772,p780,p886,p887);
FA fa228(p792,p794,p873,p888,p889);
HA ha216(p877,p881,p890,p891);
FA fa229(p883,p786,p788,p892,p893);
FA fa230(p798,p800,p802,p894,p895);
FA fa231(p804,p879,p885,p896,p897);
FA fa232(p891,p796,p810,p898,p899);
HA ha217(p887,p889,p900,p901);
HA ha218(p806,p816,p902,p903);
FA fa233(p818,p893,p895,p904,p905);
HA ha219(p897,p901,p906,p907);
FA fa234(p808,p812,p820,p908,p909);
HA ha220(p822,p899,p910,p911);
FA fa235(p903,p907,p814,p912,p913);
HA ha221(p905,p911,p914,p915);
FA fa236(p824,p830,p909,p916,p917);
HA ha222(p913,p915,p918,p919);
FA fa237(p826,p828,p834,p920,p921);
HA ha223(p836,p919,p922,p923);
HA ha224(p917,p923,p924,p925);
FA fa238(p832,p840,p921,p926,p927);
FA fa239(p925,p838,p842,p928,p929);
HA ha225(p927,p929,p930,p931);
FA fa240(p844,p931,p846,p932,p933);
FA fa241(ip_0_25,ip_1_24,ip_2_23,p934,p935);
HA ha226(ip_3_22,ip_4_21,p936,p937);
FA fa242(ip_5_20,ip_6_19,ip_7_18,p938,p939);
FA fa243(ip_8_17,ip_9_16,ip_10_15,p940,p941);
HA ha227(ip_11_14,ip_12_13,p942,p943);
FA fa244(ip_13_12,ip_14_11,ip_15_10,p944,p945);
HA ha228(ip_16_9,ip_17_8,p946,p947);
FA fa245(ip_18_7,ip_19_6,ip_20_5,p948,p949);
FA fa246(ip_21_4,ip_22_3,ip_23_2,p950,p951);
FA fa247(ip_24_1,ip_25_0,p858,p952,p953);
FA fa248(p860,p866,p937,p954,p955);
HA ha229(p943,p947,p956,p957);
HA ha230(p868,p870,p958,p959);
HA ha231(p874,p935,p960,p961);
FA fa249(p939,p941,p945,p962,p963);
HA ha232(p949,p951,p964,p965);
FA fa250(p953,p957,p850,p966,p967);
HA ha233(p852,p854,p968,p969);
HA ha234(p856,p862,p970,p971);
FA fa251(p864,p880,p882,p972,p973);
HA ha235(p955,p959,p974,p975);
FA fa252(p961,p965,p872,p976,p977);
HA ha236(p876,p890,p978,p979);
FA fa253(p963,p967,p969,p980,p981);
FA fa254(p971,p975,p878,p982,p983);
FA fa255(p884,p973,p977,p984,p985);
HA ha237(p979,p886,p986,p987);
HA ha238(p888,p900,p988,p989);
HA ha239(p981,p983,p990,p991);
HA ha240(p892,p894,p992,p993);
HA ha241(p896,p902,p994,p995);
HA ha242(p906,p985,p996,p997);
FA fa256(p987,p989,p991,p998,p999);
FA fa257(p898,p910,p993,p1000,p1001);
HA ha243(p995,p997,p1002,p1003);
HA ha244(p1003,p904,p1004,p1005);
FA fa258(p914,p999,p1001,p1006,p1007);
HA ha245(p1005,p908,p1008,p1009);
HA ha246(p912,p918,p1010,p1011);
HA ha247(p1007,p1009,p1012,p1013);
HA ha248(p1011,p922,p1014,p1015);
HA ha249(p1013,p1015,p1016,p1017);
HA ha250(p916,p924,p1018,p1019);
FA fa259(p1017,p1019,p920,p1020,p1021);
FA fa260(p1021,p926,p928,p1022,p1023);
FA fa261(p930,p1023,p932,p1024,p1025);
FA fa262(ip_0_26,ip_1_25,ip_2_24,p1026,p1027);
HA ha251(ip_3_23,ip_4_22,p1028,p1029);
HA ha252(ip_5_21,ip_6_20,p1030,p1031);
HA ha253(ip_7_19,ip_8_18,p1032,p1033);
HA ha254(ip_9_17,ip_10_16,p1034,p1035);
FA fa263(ip_11_15,ip_12_14,ip_13_13,p1036,p1037);
FA fa264(ip_14_12,ip_15_11,ip_16_10,p1038,p1039);
FA fa265(ip_17_9,ip_18_8,ip_19_7,p1040,p1041);
HA ha255(ip_20_6,ip_21_5,p1042,p1043);
FA fa266(ip_22_4,ip_23_3,ip_24_2,p1044,p1045);
HA ha256(ip_25_1,ip_26_0,p1046,p1047);
HA ha257(p1029,p1031,p1048,p1049);
FA fa267(p1033,p1035,p1043,p1050,p1051);
FA fa268(p1047,p936,p942,p1052,p1053);
HA ha258(p946,p1027,p1054,p1055);
HA ha259(p1037,p1039,p1056,p1057);
FA fa269(p1041,p1045,p1049,p1058,p1059);
FA fa270(p956,p1051,p1053,p1060,p1061);
HA ha260(p1055,p1057,p1062,p1063);
HA ha261(p934,p938,p1064,p1065);
FA fa271(p940,p944,p948,p1066,p1067);
HA ha262(p950,p952,p1068,p1069);
HA ha263(p958,p960,p1070,p1071);
FA fa272(p964,p1059,p1063,p1072,p1073);
HA ha264(p1065,p1069,p1074,p1075);
HA ha265(p1071,p954,p1076,p1077);
HA ha266(p968,p970,p1078,p1079);
FA fa273(p974,p1061,p1067,p1080,p1081);
FA fa274(p1075,p1077,p1079,p1082,p1083);
HA ha267(p962,p966,p1084,p1085);
HA ha268(p978,p1073,p1086,p1087);
HA ha269(p1085,p972,p1088,p1089);
FA fa275(p976,p1081,p1083,p1090,p1091);
HA ha270(p1087,p1089,p1092,p1093);
HA ha271(p980,p982,p1094,p1095);
FA fa276(p986,p988,p990,p1096,p1097);
HA ha272(p1093,p1095,p1098,p1099);
FA fa277(p984,p992,p994,p1100,p1101);
FA fa278(p996,p1002,p1091,p1102,p1103);
HA ha273(p1097,p1099,p1104,p1105);
HA ha274(p1004,p1101,p1106,p1107);
HA ha275(p1105,p998,p1108,p1109);
HA ha276(p1000,p1008,p1110,p1111);
HA ha277(p1010,p1103,p1112,p1113);
HA ha278(p1107,p1109,p1114,p1115);
HA ha279(p1006,p1012,p1116,p1117);
FA fa279(p1014,p1111,p1113,p1118,p1119);
HA ha280(p1115,p1016,p1120,p1121);
FA fa280(p1018,p1117,p1119,p1122,p1123);
HA ha281(p1121,p1123,p1124,p1125);
FA fa281(p1020,p1125,p1022,p1126,p1127);
HA ha282(ip_0_27,ip_1_26,p1128,p1129);
FA fa282(ip_2_25,ip_3_24,ip_4_23,p1130,p1131);
FA fa283(ip_5_22,ip_6_21,ip_7_20,p1132,p1133);
HA ha283(ip_8_19,ip_9_18,p1134,p1135);
FA fa284(ip_10_17,ip_11_16,ip_12_15,p1136,p1137);
HA ha284(ip_13_14,ip_14_13,p1138,p1139);
FA fa285(ip_15_12,ip_16_11,ip_17_10,p1140,p1141);
FA fa286(ip_18_9,ip_19_8,ip_20_7,p1142,p1143);
FA fa287(ip_21_6,ip_22_5,ip_23_4,p1144,p1145);
FA fa288(ip_24_3,ip_25_2,ip_26_1,p1146,p1147);
FA fa289(ip_27_0,p1028,p1030,p1148,p1149);
FA fa290(p1032,p1034,p1042,p1150,p1151);
HA ha285(p1046,p1129,p1152,p1153);
FA fa291(p1135,p1139,p1048,p1154,p1155);
FA fa292(p1131,p1133,p1137,p1156,p1157);
FA fa293(p1141,p1143,p1145,p1158,p1159);
FA fa294(p1147,p1153,p1026,p1160,p1161);
FA fa295(p1036,p1038,p1040,p1162,p1163);
FA fa296(p1044,p1054,p1056,p1164,p1165);
FA fa297(p1149,p1151,p1155,p1166,p1167);
FA fa298(p1050,p1052,p1062,p1168,p1169);
FA fa299(p1064,p1068,p1070,p1170,p1171);
HA ha286(p1157,p1159,p1172,p1173);
HA ha287(p1161,p1058,p1174,p1175);
HA ha288(p1074,p1076,p1176,p1177);
HA ha289(p1078,p1163,p1178,p1179);
FA fa300(p1165,p1167,p1173,p1180,p1181);
FA fa301(p1060,p1066,p1084,p1182,p1183);
HA ha290(p1169,p1171,p1184,p1185);
FA fa302(p1175,p1177,p1179,p1186,p1187);
HA ha291(p1072,p1086,p1188,p1189);
FA fa303(p1088,p1181,p1185,p1190,p1191);
FA fa304(p1080,p1082,p1092,p1192,p1193);
FA fa305(p1094,p1183,p1187,p1194,p1195);
HA ha292(p1189,p1098,p1196,p1197);
HA ha293(p1191,p1090,p1198,p1199);
HA ha294(p1096,p1104,p1200,p1201);
FA fa306(p1193,p1195,p1197,p1202,p1203);
HA ha295(p1100,p1106,p1204,p1205);
HA ha296(p1108,p1199,p1206,p1207);
HA ha297(p1201,p1102,p1208,p1209);
FA fa307(p1110,p1112,p1114,p1210,p1211);
FA fa308(p1203,p1205,p1207,p1212,p1213);
HA ha298(p1116,p1209,p1214,p1215);
HA ha299(p1120,p1211,p1216,p1217);
FA fa309(p1213,p1215,p1118,p1218,p1219);
HA ha300(p1217,p1122,p1220,p1221);
HA ha301(p1124,p1219,p1222,p1223);
HA ha302(p1221,p1223,p1224,p1225);
FA fa310(ip_0_28,ip_1_27,ip_2_26,p1226,p1227);
HA ha303(ip_3_25,ip_4_24,p1228,p1229);
FA fa311(ip_5_23,ip_6_22,ip_7_21,p1230,p1231);
FA fa312(ip_8_20,ip_9_19,ip_10_18,p1232,p1233);
HA ha304(ip_11_17,ip_12_16,p1234,p1235);
HA ha305(ip_13_15,ip_14_14,p1236,p1237);
HA ha306(ip_15_13,ip_16_12,p1238,p1239);
HA ha307(ip_17_11,ip_18_10,p1240,p1241);
FA fa313(ip_19_9,ip_20_8,ip_21_7,p1242,p1243);
HA ha308(ip_22_6,ip_23_5,p1244,p1245);
HA ha309(ip_24_4,ip_25_3,p1246,p1247);
HA ha310(ip_26_2,ip_27_1,p1248,p1249);
FA fa314(ip_28_0,p1128,p1134,p1250,p1251);
FA fa315(p1138,p1229,p1235,p1252,p1253);
HA ha311(p1237,p1239,p1254,p1255);
HA ha312(p1241,p1245,p1256,p1257);
FA fa316(p1247,p1249,p1152,p1258,p1259);
FA fa317(p1227,p1231,p1233,p1260,p1261);
FA fa318(p1243,p1255,p1257,p1262,p1263);
FA fa319(p1130,p1132,p1136,p1264,p1265);
HA ha313(p1140,p1142,p1266,p1267);
FA fa320(p1144,p1146,p1251,p1268,p1269);
HA ha314(p1253,p1259,p1270,p1271);
HA ha315(p1148,p1150,p1272,p1273);
HA ha316(p1154,p1261,p1274,p1275);
FA fa321(p1263,p1267,p1271,p1276,p1277);
FA fa322(p1156,p1158,p1160,p1278,p1279);
HA ha317(p1172,p1265,p1280,p1281);
HA ha318(p1269,p1273,p1282,p1283);
FA fa323(p1275,p1162,p1164,p1284,p1285);
FA fa324(p1166,p1174,p1176,p1286,p1287);
HA ha319(p1178,p1277,p1288,p1289);
HA ha320(p1281,p1283,p1290,p1291);
FA fa325(p1168,p1170,p1184,p1292,p1293);
FA fa326(p1279,p1289,p1291,p1294,p1295);
HA ha321(p1180,p1188,p1296,p1297);
FA fa327(p1285,p1287,p1182,p1298,p1299);
FA fa328(p1186,p1293,p1295,p1300,p1301);
FA fa329(p1297,p1190,p1196,p1302,p1303);
HA ha322(p1299,p1192,p1304,p1305);
HA ha323(p1194,p1198,p1306,p1307);
HA ha324(p1200,p1301,p1308,p1309);
HA ha325(p1204,p1206,p1310,p1311);
HA ha326(p1303,p1305,p1312,p1313);
FA fa330(p1307,p1309,p1202,p1314,p1315);
FA fa331(p1208,p1311,p1313,p1316,p1317);
FA fa332(p1214,p1315,p1210,p1318,p1319);
HA ha327(p1212,p1216,p1320,p1321);
HA ha328(p1317,p1319,p1322,p1323);
HA ha329(p1321,p1218,p1324,p1325);
HA ha330(p1220,p1222,p1326,p1327);
HA ha331(p1323,p1224,p1328,p1329);
HA ha332(p1325,p1327,p1330,p1331);
HA ha333(ip_0_29,ip_1_28,p1332,p1333);
HA ha334(ip_2_27,ip_3_26,p1334,p1335);
HA ha335(ip_4_25,ip_5_24,p1336,p1337);
HA ha336(ip_6_23,ip_7_22,p1338,p1339);
HA ha337(ip_8_21,ip_9_20,p1340,p1341);
FA fa333(ip_10_19,ip_11_18,ip_12_17,p1342,p1343);
HA ha338(ip_13_16,ip_14_15,p1344,p1345);
HA ha339(ip_15_14,ip_16_13,p1346,p1347);
HA ha340(ip_17_12,ip_18_11,p1348,p1349);
FA fa334(ip_19_10,ip_20_9,ip_21_8,p1350,p1351);
HA ha341(ip_22_7,ip_23_6,p1352,p1353);
HA ha342(ip_24_5,ip_25_4,p1354,p1355);
HA ha343(ip_26_3,ip_27_2,p1356,p1357);
HA ha344(ip_28_1,ip_29_0,p1358,p1359);
HA ha345(p1228,p1234,p1360,p1361);
HA ha346(p1236,p1238,p1362,p1363);
FA fa335(p1240,p1244,p1246,p1364,p1365);
HA ha347(p1248,p1333,p1366,p1367);
HA ha348(p1335,p1337,p1368,p1369);
HA ha349(p1339,p1341,p1370,p1371);
FA fa336(p1345,p1347,p1349,p1372,p1373);
FA fa337(p1353,p1355,p1357,p1374,p1375);
HA ha350(p1359,p1254,p1376,p1377);
HA ha351(p1256,p1343,p1378,p1379);
FA fa338(p1351,p1361,p1363,p1380,p1381);
HA ha352(p1367,p1369,p1382,p1383);
HA ha353(p1371,p1226,p1384,p1385);
HA ha354(p1230,p1232,p1386,p1387);
FA fa339(p1242,p1365,p1373,p1388,p1389);
HA ha355(p1375,p1377,p1390,p1391);
HA ha356(p1379,p1383,p1392,p1393);
FA fa340(p1250,p1252,p1258,p1394,p1395);
HA ha357(p1266,p1270,p1396,p1397);
FA fa341(p1381,p1385,p1387,p1398,p1399);
FA fa342(p1391,p1393,p1260,p1400,p1401);
HA ha358(p1262,p1272,p1402,p1403);
HA ha359(p1274,p1389,p1404,p1405);
FA fa343(p1397,p1264,p1268,p1406,p1407);
FA fa344(p1280,p1282,p1395,p1408,p1409);
HA ha360(p1399,p1401,p1410,p1411);
FA fa345(p1403,p1405,p1276,p1412,p1413);
HA ha361(p1288,p1290,p1414,p1415);
HA ha362(p1411,p1278,p1416,p1417);
HA ha363(p1407,p1409,p1418,p1419);
FA fa346(p1413,p1415,p1284,p1420,p1421);
HA ha364(p1286,p1296,p1422,p1423);
HA ha365(p1417,p1419,p1424,p1425);
FA fa347(p1292,p1294,p1421,p1426,p1427);
HA ha366(p1423,p1425,p1428,p1429);
FA fa348(p1298,p1429,p1300,p1430,p1431);
HA ha367(p1304,p1306,p1432,p1433);
HA ha368(p1308,p1427,p1434,p1435);
HA ha369(p1302,p1310,p1436,p1437);
HA ha370(p1312,p1431,p1438,p1439);
HA ha371(p1433,p1435,p1440,p1441);
FA fa349(p1437,p1439,p1441,p1442,p1443);
HA ha372(p1314,p1316,p1444,p1445);
HA ha373(p1320,p1443,p1446,p1447);
FA fa350(p1318,p1322,p1445,p1448,p1449);
FA fa351(p1447,p1324,p1326,p1450,p1451);
FA fa352(p1328,p1330,p1449,p1452,p1453);
FA fa353(ip_0_30,ip_1_29,ip_2_28,p1454,p1455);
HA ha374(ip_3_27,ip_4_26,p1456,p1457);
FA fa354(ip_5_25,ip_6_24,ip_7_23,p1458,p1459);
FA fa355(ip_8_22,ip_9_21,ip_10_20,p1460,p1461);
FA fa356(ip_11_19,ip_12_18,ip_13_17,p1462,p1463);
FA fa357(ip_14_16,ip_15_15,ip_16_14,p1464,p1465);
HA ha375(ip_17_13,ip_18_12,p1466,p1467);
HA ha376(ip_19_11,ip_20_10,p1468,p1469);
HA ha377(ip_21_9,ip_22_8,p1470,p1471);
HA ha378(ip_23_7,ip_24_6,p1472,p1473);
HA ha379(ip_25_5,ip_26_4,p1474,p1475);
HA ha380(ip_27_3,ip_28_2,p1476,p1477);
HA ha381(ip_29_1,ip_30_0,p1478,p1479);
FA fa358(p1332,p1334,p1336,p1480,p1481);
FA fa359(p1338,p1340,p1344,p1482,p1483);
FA fa360(p1346,p1348,p1352,p1484,p1485);
HA ha382(p1354,p1356,p1486,p1487);
HA ha383(p1358,p1457,p1488,p1489);
HA ha384(p1467,p1469,p1490,p1491);
HA ha385(p1471,p1473,p1492,p1493);
HA ha386(p1475,p1477,p1494,p1495);
HA ha387(p1479,p1360,p1496,p1497);
FA fa361(p1362,p1366,p1368,p1498,p1499);
HA ha388(p1370,p1455,p1500,p1501);
HA ha389(p1459,p1461,p1502,p1503);
FA fa362(p1463,p1465,p1487,p1504,p1505);
HA ha390(p1489,p1491,p1506,p1507);
FA fa363(p1493,p1495,p1342,p1508,p1509);
HA ha391(p1350,p1376,p1510,p1511);
FA fa364(p1378,p1382,p1481,p1512,p1513);
FA fa365(p1483,p1485,p1497,p1514,p1515);
HA ha392(p1501,p1503,p1516,p1517);
FA fa366(p1507,p1364,p1372,p1518,p1519);
FA fa367(p1374,p1384,p1386,p1520,p1521);
HA ha393(p1390,p1392,p1522,p1523);
HA ha394(p1499,p1505,p1524,p1525);
HA ha395(p1509,p1511,p1526,p1527);
HA ha396(p1517,p1380,p1528,p1529);
HA ha397(p1396,p1513,p1530,p1531);
FA fa368(p1515,p1523,p1525,p1532,p1533);
FA fa369(p1527,p1388,p1402,p1534,p1535);
HA ha398(p1404,p1519,p1536,p1537);
FA fa370(p1521,p1529,p1531,p1538,p1539);
HA ha399(p1394,p1398,p1540,p1541);
HA ha400(p1400,p1410,p1542,p1543);
HA ha401(p1533,p1537,p1544,p1545);
HA ha402(p1414,p1535,p1546,p1547);
FA fa371(p1539,p1541,p1543,p1548,p1549);
HA ha403(p1545,p1406,p1550,p1551);
HA ha404(p1408,p1412,p1552,p1553);
FA fa372(p1416,p1418,p1547,p1554,p1555);
FA fa373(p1422,p1424,p1549,p1556,p1557);
HA ha405(p1551,p1553,p1558,p1559);
HA ha406(p1420,p1428,p1560,p1561);
FA fa374(p1555,p1559,p1557,p1562,p1563);
HA ha407(p1561,p1426,p1564,p1565);
HA ha408(p1432,p1434,p1566,p1567);
HA ha409(p1563,p1430,p1568,p1569);
HA ha410(p1436,p1438,p1570,p1571);
HA ha411(p1440,p1565,p1572,p1573);
HA ha412(p1567,p1569,p1574,p1575);
FA fa375(p1571,p1573,p1575,p1576,p1577);
HA ha413(p1442,p1444,p1578,p1579);
FA fa376(p1446,p1577,p1579,p1580,p1581);
FA fa377(p1581,p1448,p1450,p1582,p1583);
HA ha414(ip_0_31,ip_1_30,p1584,p1585);
HA ha415(ip_2_29,ip_3_28,p1586,p1587);
FA fa378(ip_4_27,ip_5_26,ip_6_25,p1588,p1589);
FA fa379(ip_7_24,ip_8_23,ip_9_22,p1590,p1591);
HA ha416(ip_10_21,ip_11_20,p1592,p1593);
FA fa380(ip_12_19,ip_13_18,ip_14_17,p1594,p1595);
FA fa381(ip_15_16,ip_16_15,ip_17_14,p1596,p1597);
HA ha417(ip_18_13,ip_19_12,p1598,p1599);
HA ha418(ip_20_11,ip_21_10,p1600,p1601);
HA ha419(ip_22_9,ip_23_8,p1602,p1603);
HA ha420(ip_24_7,ip_25_6,p1604,p1605);
FA fa382(ip_26_5,ip_27_4,ip_28_3,p1606,p1607);
FA fa383(ip_29_2,ip_30_1,ip_31_0,p1608,p1609);
HA ha421(p1456,p1466,p1610,p1611);
FA fa384(p1468,p1470,p1472,p1612,p1613);
FA fa385(p1474,p1476,p1478,p1614,p1615);
HA ha422(p1585,p1587,p1616,p1617);
HA ha423(p1593,p1599,p1618,p1619);
FA fa386(p1601,p1603,p1605,p1620,p1621);
HA ha424(p1486,p1488,p1622,p1623);
HA ha425(p1490,p1492,p1624,p1625);
FA fa387(p1494,p1589,p1591,p1626,p1627);
FA fa388(p1595,p1597,p1607,p1628,p1629);
FA fa389(p1609,p1611,p1617,p1630,p1631);
FA fa390(p1619,p1454,p1458,p1632,p1633);
FA fa391(p1460,p1462,p1464,p1634,p1635);
FA fa392(p1496,p1500,p1502,p1636,p1637);
HA ha426(p1506,p1613,p1638,p1639);
HA ha427(p1615,p1621,p1640,p1641);
FA fa393(p1623,p1625,p1480,p1642,p1643);
FA fa394(p1482,p1484,p1510,p1644,p1645);
FA fa395(p1516,p1627,p1629,p1646,p1647);
HA ha428(p1631,p1639,p1648,p1649);
HA ha429(p1641,p1498,p1650,p1651);
FA fa396(p1504,p1508,p1522,p1652,p1653);
FA fa397(p1524,p1526,p1633,p1654,p1655);
HA ha430(p1635,p1637,p1656,p1657);
HA ha431(p1643,p1649,p1658,p1659);
FA fa398(p1512,p1514,p1528,p1660,p1661);
FA fa399(p1530,p1645,p1647,p1662,p1663);
HA ha432(p1651,p1657,p1664,p1665);
HA ha433(p1659,p1518,p1666,p1667);
HA ha434(p1520,p1536,p1668,p1669);
FA fa400(p1653,p1655,p1665,p1670,p1671);
HA ha435(p1532,p1540,p1672,p1673);
FA fa401(p1542,p1544,p1661,p1674,p1675);
HA ha436(p1663,p1667,p1676,p1677);
HA ha437(p1669,p1534,p1678,p1679);
FA fa402(p1538,p1546,p1671,p1680,p1681);
FA fa403(p1673,p1677,p1550,p1682,p1683);
HA ha438(p1552,p1675,p1684,p1685);
HA ha439(p1679,p1548,p1686,p1687);
HA ha440(p1558,p1681,p1688,p1689);
HA ha441(p1683,p1685,p1690,p1691);
FA fa404(p1554,p1560,p1687,p1692,p1693);
FA fa405(p1689,p1691,p1556,p1694,p1695);
FA fa406(p1562,p1564,p1566,p1696,p1697);
FA fa407(p1693,p1695,p1568,p1698,p1699);
HA ha442(p1570,p1572,p1700,p1701);
HA ha443(p1574,p1697,p1702,p1703);
FA fa408(p1699,p1701,p1703,p1704,p1705);
HA ha444(p1576,p1578,p1706,p1707);
HA ha445(p1705,p1707,p1708,p1709);
FA fa409(p1580,p1709,p1582,p1710,p1711);
HA ha446(ip_1_31,ip_2_30,p1712,p1713);
FA fa410(ip_3_29,ip_4_28,ip_5_27,p1714,p1715);
FA fa411(ip_6_26,ip_7_25,ip_8_24,p1716,p1717);
FA fa412(ip_9_23,ip_10_22,ip_11_21,p1718,p1719);
FA fa413(ip_12_20,ip_13_19,ip_14_18,p1720,p1721);
HA ha447(ip_15_17,ip_16_16,p1722,p1723);
FA fa414(ip_17_15,ip_18_14,ip_19_13,p1724,p1725);
HA ha448(ip_20_12,ip_21_11,p1726,p1727);
HA ha449(ip_22_10,ip_23_9,p1728,p1729);
HA ha450(ip_24_8,ip_25_7,p1730,p1731);
FA fa415(ip_26_6,ip_27_5,ip_28_4,p1732,p1733);
HA ha451(ip_29_3,ip_30_2,p1734,p1735);
FA fa416(ip_31_1,p1584,p1586,p1736,p1737);
HA ha452(p1592,p1598,p1738,p1739);
HA ha453(p1600,p1602,p1740,p1741);
FA fa417(p1604,p1713,p1723,p1742,p1743);
FA fa418(p1727,p1729,p1731,p1744,p1745);
HA ha454(p1735,p1610,p1746,p1747);
HA ha455(p1616,p1618,p1748,p1749);
HA ha456(p1715,p1717,p1750,p1751);
FA fa419(p1719,p1721,p1725,p1752,p1753);
HA ha457(p1733,p1739,p1754,p1755);
HA ha458(p1741,p1588,p1756,p1757);
HA ha459(p1590,p1594,p1758,p1759);
FA fa420(p1596,p1606,p1608,p1760,p1761);
HA ha460(p1622,p1624,p1762,p1763);
FA fa421(p1737,p1743,p1745,p1764,p1765);
FA fa422(p1747,p1749,p1751,p1766,p1767);
FA fa423(p1755,p1612,p1614,p1768,p1769);
HA ha461(p1620,p1638,p1770,p1771);
FA fa424(p1640,p1753,p1757,p1772,p1773);
HA ha462(p1759,p1763,p1774,p1775);
HA ha463(p1626,p1628,p1776,p1777);
HA ha464(p1630,p1648,p1778,p1779);
HA ha465(p1761,p1765,p1780,p1781);
FA fa425(p1767,p1771,p1775,p1782,p1783);
HA ha466(p1632,p1634,p1784,p1785);
HA ha467(p1636,p1642,p1786,p1787);
FA fa426(p1650,p1656,p1658,p1788,p1789);
HA ha468(p1769,p1773,p1790,p1791);
FA fa427(p1777,p1779,p1781,p1792,p1793);
FA fa428(p1644,p1646,p1664,p1794,p1795);
HA ha469(p1783,p1785,p1796,p1797);
HA ha470(p1787,p1791,p1798,p1799);
FA fa429(p1652,p1654,p1666,p1800,p1801);
HA ha471(p1668,p1789,p1802,p1803);
FA fa430(p1793,p1797,p1799,p1804,p1805);
FA fa431(p1660,p1662,p1672,p1806,p1807);
FA fa432(p1676,p1795,p1803,p1808,p1809);
FA fa433(p1670,p1678,p1801,p1810,p1811);
FA fa434(p1805,p1674,p1684,p1812,p1813);
HA ha472(p1807,p1809,p1814,p1815);
FA fa435(p1680,p1682,p1686,p1816,p1817);
HA ha473(p1688,p1690,p1818,p1819);
FA fa436(p1811,p1815,p1813,p1820,p1821);
HA ha474(p1819,p1817,p1822,p1823);
HA ha475(p1821,p1692,p1824,p1825);
HA ha476(p1694,p1823,p1826,p1827);
HA ha477(p1700,p1825,p1828,p1829);
HA ha478(p1827,p1696,p1830,p1831);
HA ha479(p1698,p1702,p1832,p1833);
HA ha480(p1829,p1831,p1834,p1835);
HA ha481(p1833,p1704,p1836,p1837);
HA ha482(p1706,p1835,p1838,p1839);
FA fa437(p1708,p1837,p1839,p1840,p1841);
HA ha483(ip_2_31,ip_3_30,p1842,p1843);
FA fa438(ip_4_29,ip_5_28,ip_6_27,p1844,p1845);
FA fa439(ip_7_26,ip_8_25,ip_9_24,p1846,p1847);
HA ha484(ip_10_23,ip_11_22,p1848,p1849);
FA fa440(ip_12_21,ip_13_20,ip_14_19,p1850,p1851);
FA fa441(ip_15_18,ip_16_17,ip_17_16,p1852,p1853);
HA ha485(ip_18_15,ip_19_14,p1854,p1855);
FA fa442(ip_20_13,ip_21_12,ip_22_11,p1856,p1857);
FA fa443(ip_23_10,ip_24_9,ip_25_8,p1858,p1859);
HA ha486(ip_26_7,ip_27_6,p1860,p1861);
FA fa444(ip_28_5,ip_29_4,ip_30_3,p1862,p1863);
FA fa445(ip_31_2,p1712,p1722,p1864,p1865);
HA ha487(p1726,p1728,p1866,p1867);
FA fa446(p1730,p1734,p1843,p1868,p1869);
HA ha488(p1849,p1855,p1870,p1871);
FA fa447(p1861,p1738,p1740,p1872,p1873);
HA ha489(p1845,p1847,p1874,p1875);
HA ha490(p1851,p1853,p1876,p1877);
FA fa448(p1857,p1859,p1863,p1878,p1879);
FA fa449(p1867,p1871,p1714,p1880,p1881);
HA ha491(p1716,p1718,p1882,p1883);
HA ha492(p1720,p1724,p1884,p1885);
FA fa450(p1732,p1746,p1748,p1886,p1887);
HA ha493(p1750,p1754,p1888,p1889);
HA ha494(p1865,p1869,p1890,p1891);
FA fa451(p1875,p1877,p1736,p1892,p1893);
HA ha495(p1742,p1744,p1894,p1895);
HA ha496(p1756,p1758,p1896,p1897);
HA ha497(p1762,p1873,p1898,p1899);
HA ha498(p1879,p1881,p1900,p1901);
FA fa452(p1883,p1885,p1889,p1902,p1903);
HA ha499(p1891,p1752,p1904,p1905);
FA fa453(p1770,p1774,p1887,p1906,p1907);
FA fa454(p1893,p1895,p1897,p1908,p1909);
HA ha500(p1899,p1901,p1910,p1911);
HA ha501(p1760,p1764,p1912,p1913);
HA ha502(p1766,p1776,p1914,p1915);
HA ha503(p1778,p1780,p1916,p1917);
HA ha504(p1903,p1905,p1918,p1919);
HA ha505(p1911,p1768,p1920,p1921);
HA ha506(p1772,p1784,p1922,p1923);
HA ha507(p1786,p1790,p1924,p1925);
FA fa455(p1907,p1909,p1913,p1926,p1927);
HA ha508(p1915,p1917,p1928,p1929);
HA ha509(p1919,p1782,p1930,p1931);
HA ha510(p1796,p1798,p1932,p1933);
HA ha511(p1921,p1923,p1934,p1935);
HA ha512(p1925,p1929,p1936,p1937);
HA ha513(p1788,p1792,p1938,p1939);
FA fa456(p1802,p1927,p1931,p1940,p1941);
FA fa457(p1933,p1935,p1937,p1942,p1943);
FA fa458(p1794,p1939,p1800,p1944,p1945);
HA ha514(p1804,p1941,p1946,p1947);
FA fa459(p1943,p1806,p1808,p1948,p1949);
HA ha515(p1814,p1945,p1950,p1951);
FA fa460(p1947,p1810,p1818,p1952,p1953);
HA ha516(p1951,p1812,p1954,p1955);
HA ha517(p1949,p1816,p1956,p1957);
HA ha518(p1820,p1822,p1958,p1959);
HA ha519(p1953,p1955,p1960,p1961);
HA ha520(p1824,p1826,p1962,p1963);
HA ha521(p1957,p1959,p1964,p1965);
FA fa461(p1961,p1828,p1963,p1966,p1967);
HA ha522(p1965,p1830,p1968,p1969);
HA ha523(p1832,p1834,p1970,p1971);
FA fa462(p1967,p1969,p1836,p1972,p1973);
FA fa463(p1838,p1971,p1973,p1974,p1975);
FA fa464(ip_3_31,ip_4_30,ip_5_29,p1976,p1977);
HA ha524(ip_6_28,ip_7_27,p1978,p1979);
HA ha525(ip_8_26,ip_9_25,p1980,p1981);
HA ha526(ip_10_24,ip_11_23,p1982,p1983);
HA ha527(ip_12_22,ip_13_21,p1984,p1985);
FA fa465(ip_14_20,ip_15_19,ip_16_18,p1986,p1987);
HA ha528(ip_17_17,ip_18_16,p1988,p1989);
HA ha529(ip_19_15,ip_20_14,p1990,p1991);
HA ha530(ip_21_13,ip_22_12,p1992,p1993);
FA fa466(ip_23_11,ip_24_10,ip_25_9,p1994,p1995);
FA fa467(ip_26_8,ip_27_7,ip_28_6,p1996,p1997);
FA fa468(ip_29_5,ip_30_4,ip_31_3,p1998,p1999);
HA ha531(p1842,p1848,p2000,p2001);
FA fa469(p1854,p1860,p1979,p2002,p2003);
FA fa470(p1981,p1983,p1985,p2004,p2005);
FA fa471(p1989,p1991,p1993,p2006,p2007);
HA ha532(p1866,p1870,p2008,p2009);
FA fa472(p1977,p1987,p1995,p2010,p2011);
HA ha533(p1997,p1999,p2012,p2013);
FA fa473(p2001,p1844,p1846,p2014,p2015);
FA fa474(p1850,p1852,p1856,p2016,p2017);
FA fa475(p1858,p1862,p1874,p2018,p2019);
FA fa476(p1876,p2003,p2005,p2020,p2021);
HA ha534(p2007,p2009,p2022,p2023);
HA ha535(p2013,p1864,p2024,p2025);
FA fa477(p1868,p1882,p1884,p2026,p2027);
HA ha536(p1888,p1890,p2028,p2029);
HA ha537(p2011,p2023,p2030,p2031);
HA ha538(p1872,p1878,p2032,p2033);
FA fa478(p1880,p1894,p1896,p2034,p2035);
HA ha539(p1898,p1900,p2036,p2037);
FA fa479(p2015,p2017,p2019,p2038,p2039);
FA fa480(p2021,p2025,p2029,p2040,p2041);
HA ha540(p2031,p1886,p2042,p2043);
HA ha541(p1892,p1904,p2044,p2045);
FA fa481(p1910,p2027,p2033,p2046,p2047);
HA ha542(p2037,p1902,p2048,p2049);
FA fa482(p1912,p1914,p1916,p2050,p2051);
HA ha543(p1918,p2035,p2052,p2053);
HA ha544(p2039,p2041,p2054,p2055);
FA fa483(p2043,p2045,p1906,p2056,p2057);
HA ha545(p1908,p1920,p2058,p2059);
FA fa484(p1922,p1924,p1928,p2060,p2061);
HA ha546(p2047,p2049,p2062,p2063);
HA ha547(p2053,p2055,p2064,p2065);
HA ha548(p1930,p1932,p2066,p2067);
HA ha549(p1934,p1936,p2068,p2069);
HA ha550(p2051,p2057,p2070,p2071);
HA ha551(p2059,p2063,p2072,p2073);
HA ha552(p2065,p1926,p2074,p2075);
HA ha553(p1938,p2061,p2076,p2077);
FA fa485(p2067,p2069,p2071,p2078,p2079);
FA fa486(p2073,p2075,p2077,p2080,p2081);
HA ha554(p1940,p1942,p2082,p2083);
HA ha555(p1946,p2079,p2084,p2085);
HA ha556(p1944,p1950,p2086,p2087);
FA fa487(p2081,p2083,p2085,p2088,p2089);
FA fa488(p2087,p1948,p1954,p2090,p2091);
HA ha557(p2089,p1952,p2092,p2093);
FA fa489(p1956,p1958,p1960,p2094,p2095);
HA ha558(p1962,p1964,p2096,p2097);
FA fa490(p2091,p2093,p2095,p2098,p2099);
HA ha559(p2097,p1968,p2100,p2101);
FA fa491(p2099,p1966,p1970,p2102,p2103);
HA ha560(p2101,p1972,p2104,p2105);
FA fa492(p2103,p1974,p2105,p2106,p2107);
FA fa493(ip_4_31,ip_5_30,ip_6_29,p2108,p2109);
HA ha561(ip_7_28,ip_8_27,p2110,p2111);
FA fa494(ip_9_26,ip_10_25,ip_11_24,p2112,p2113);
HA ha562(ip_12_23,ip_13_22,p2114,p2115);
HA ha563(ip_14_21,ip_15_20,p2116,p2117);
HA ha564(ip_16_19,ip_17_18,p2118,p2119);
FA fa495(ip_18_17,ip_19_16,ip_20_15,p2120,p2121);
HA ha565(ip_21_14,ip_22_13,p2122,p2123);
HA ha566(ip_23_12,ip_24_11,p2124,p2125);
FA fa496(ip_25_10,ip_26_9,ip_27_8,p2126,p2127);
HA ha567(ip_28_7,ip_29_6,p2128,p2129);
HA ha568(ip_30_5,ip_31_4,p2130,p2131);
FA fa497(p1978,p1980,p1982,p2132,p2133);
HA ha569(p1984,p1988,p2134,p2135);
HA ha570(p1990,p1992,p2136,p2137);
HA ha571(p2111,p2115,p2138,p2139);
HA ha572(p2117,p2119,p2140,p2141);
HA ha573(p2123,p2125,p2142,p2143);
HA ha574(p2129,p2131,p2144,p2145);
HA ha575(p2000,p2109,p2146,p2147);
FA fa498(p2113,p2121,p2127,p2148,p2149);
HA ha576(p2135,p2137,p2150,p2151);
HA ha577(p2139,p2141,p2152,p2153);
FA fa499(p2143,p2145,p1976,p2154,p2155);
HA ha578(p1986,p1994,p2156,p2157);
HA ha579(p1996,p1998,p2158,p2159);
FA fa500(p2008,p2012,p2133,p2160,p2161);
HA ha580(p2147,p2151,p2162,p2163);
HA ha581(p2153,p2002,p2164,p2165);
HA ha582(p2004,p2006,p2166,p2167);
FA fa501(p2022,p2149,p2155,p2168,p2169);
HA ha583(p2157,p2159,p2170,p2171);
HA ha584(p2163,p2010,p2172,p2173);
HA ha585(p2024,p2028,p2174,p2175);
FA fa502(p2030,p2161,p2165,p2176,p2177);
HA ha586(p2167,p2171,p2178,p2179);
FA fa503(p2014,p2016,p2018,p2180,p2181);
FA fa504(p2020,p2032,p2036,p2182,p2183);
FA fa505(p2169,p2173,p2175,p2184,p2185);
HA ha587(p2179,p2026,p2186,p2187);
HA ha588(p2042,p2044,p2188,p2189);
HA ha589(p2177,p2034,p2190,p2191);
FA fa506(p2038,p2040,p2048,p2192,p2193);
HA ha590(p2052,p2054,p2194,p2195);
HA ha591(p2181,p2183,p2196,p2197);
HA ha592(p2185,p2187,p2198,p2199);
HA ha593(p2189,p2046,p2200,p2201);
FA fa507(p2058,p2062,p2064,p2202,p2203);
FA fa508(p2191,p2195,p2197,p2204,p2205);
FA fa509(p2199,p2050,p2056,p2206,p2207);
FA fa510(p2066,p2068,p2070,p2208,p2209);
HA ha594(p2072,p2193,p2210,p2211);
HA ha595(p2201,p2060,p2212,p2213);
FA fa511(p2074,p2076,p2203,p2214,p2215);
FA fa512(p2205,p2211,p2207,p2216,p2217);
FA fa513(p2209,p2213,p2078,p2218,p2219);
FA fa514(p2082,p2084,p2215,p2220,p2221);
FA fa515(p2217,p2080,p2086,p2222,p2223);
FA fa516(p2219,p2221,p2088,p2224,p2225);
HA ha596(p2223,p2092,p2226,p2227);
FA fa517(p2225,p2090,p2096,p2228,p2229);
HA ha597(p2227,p2094,p2230,p2231);
HA ha598(p2098,p2100,p2232,p2233);
FA fa518(p2229,p2231,p2233,p2234,p2235);
HA ha599(p2235,p2102,p2236,p2237);
HA ha600(p2104,p2237,p2238,p2239);
HA ha601(ip_5_31,ip_6_30,p2240,p2241);
HA ha602(ip_7_29,ip_8_28,p2242,p2243);
FA fa519(ip_9_27,ip_10_26,ip_11_25,p2244,p2245);
FA fa520(ip_12_24,ip_13_23,ip_14_22,p2246,p2247);
HA ha603(ip_15_21,ip_16_20,p2248,p2249);
FA fa521(ip_17_19,ip_18_18,ip_19_17,p2250,p2251);
HA ha604(ip_20_16,ip_21_15,p2252,p2253);
FA fa522(ip_22_14,ip_23_13,ip_24_12,p2254,p2255);
FA fa523(ip_25_11,ip_26_10,ip_27_9,p2256,p2257);
HA ha605(ip_28_8,ip_29_7,p2258,p2259);
FA fa524(ip_30_6,ip_31_5,p2110,p2260,p2261);
HA ha606(p2114,p2116,p2262,p2263);
HA ha607(p2118,p2122,p2264,p2265);
HA ha608(p2124,p2128,p2266,p2267);
HA ha609(p2130,p2241,p2268,p2269);
HA ha610(p2243,p2249,p2270,p2271);
HA ha611(p2253,p2259,p2272,p2273);
FA fa525(p2134,p2136,p2138,p2274,p2275);
FA fa526(p2140,p2142,p2144,p2276,p2277);
HA ha612(p2245,p2247,p2278,p2279);
HA ha613(p2251,p2255,p2280,p2281);
HA ha614(p2257,p2261,p2282,p2283);
FA fa527(p2263,p2265,p2267,p2284,p2285);
HA ha615(p2269,p2271,p2286,p2287);
HA ha616(p2273,p2108,p2288,p2289);
FA fa528(p2112,p2120,p2126,p2290,p2291);
FA fa529(p2146,p2150,p2152,p2292,p2293);
HA ha617(p2279,p2281,p2294,p2295);
HA ha618(p2283,p2287,p2296,p2297);
FA fa530(p2132,p2156,p2158,p2298,p2299);
FA fa531(p2162,p2275,p2277,p2300,p2301);
HA ha619(p2285,p2289,p2302,p2303);
HA ha620(p2295,p2297,p2304,p2305);
HA ha621(p2148,p2154,p2306,p2307);
FA fa532(p2164,p2166,p2170,p2308,p2309);
FA fa533(p2291,p2293,p2303,p2310,p2311);
FA fa534(p2305,p2160,p2172,p2312,p2313);
HA ha622(p2174,p2178,p2314,p2315);
FA fa535(p2299,p2301,p2307,p2316,p2317);
FA fa536(p2168,p2309,p2311,p2318,p2319);
FA fa537(p2315,p2176,p2186,p2320,p2321);
FA fa538(p2188,p2313,p2317,p2322,p2323);
FA fa539(p2180,p2182,p2184,p2324,p2325);
FA fa540(p2190,p2194,p2196,p2326,p2327);
FA fa541(p2198,p2319,p2200,p2328,p2329);
HA ha623(p2321,p2323,p2330,p2331);
FA fa542(p2192,p2210,p2325,p2332,p2333);
FA fa543(p2327,p2329,p2331,p2334,p2335);
HA ha624(p2202,p2204,p2336,p2337);
FA fa544(p2212,p2206,p2208,p2338,p2339);
FA fa545(p2333,p2335,p2337,p2340,p2341);
FA fa546(p2214,p2216,p2218,p2342,p2343);
HA ha625(p2339,p2341,p2344,p2345);
HA ha626(p2220,p2343,p2346,p2347);
FA fa547(p2345,p2222,p2347,p2348,p2349);
FA fa548(p2224,p2226,p2349,p2350,p2351);
HA ha627(p2230,p2351,p2352,p2353);
FA fa549(p2228,p2232,p2353,p2354,p2355);
FA fa550(p2234,p2355,p2236,p2356,p2357);
HA ha628(ip_6_31,ip_7_30,p2358,p2359);
HA ha629(ip_8_29,ip_9_28,p2360,p2361);
HA ha630(ip_10_27,ip_11_26,p2362,p2363);
HA ha631(ip_12_25,ip_13_24,p2364,p2365);
HA ha632(ip_14_23,ip_15_22,p2366,p2367);
HA ha633(ip_16_21,ip_17_20,p2368,p2369);
HA ha634(ip_18_19,ip_19_18,p2370,p2371);
HA ha635(ip_20_17,ip_21_16,p2372,p2373);
HA ha636(ip_22_15,ip_23_14,p2374,p2375);
HA ha637(ip_24_13,ip_25_12,p2376,p2377);
HA ha638(ip_26_11,ip_27_10,p2378,p2379);
HA ha639(ip_28_9,ip_29_8,p2380,p2381);
FA fa551(ip_30_7,ip_31_6,p2240,p2382,p2383);
HA ha640(p2242,p2248,p2384,p2385);
HA ha641(p2252,p2258,p2386,p2387);
HA ha642(p2359,p2361,p2388,p2389);
HA ha643(p2363,p2365,p2390,p2391);
HA ha644(p2367,p2369,p2392,p2393);
FA fa552(p2371,p2373,p2375,p2394,p2395);
FA fa553(p2377,p2379,p2381,p2396,p2397);
FA fa554(p2262,p2264,p2266,p2398,p2399);
HA ha645(p2268,p2270,p2400,p2401);
FA fa555(p2272,p2383,p2385,p2402,p2403);
FA fa556(p2387,p2389,p2391,p2404,p2405);
FA fa557(p2393,p2244,p2246,p2406,p2407);
FA fa558(p2250,p2254,p2256,p2408,p2409);
FA fa559(p2260,p2278,p2280,p2410,p2411);
HA ha646(p2282,p2286,p2412,p2413);
HA ha647(p2395,p2397,p2414,p2415);
HA ha648(p2401,p2288,p2416,p2417);
HA ha649(p2294,p2296,p2418,p2419);
FA fa560(p2399,p2403,p2405,p2420,p2421);
HA ha650(p2413,p2415,p2422,p2423);
FA fa561(p2274,p2276,p2284,p2424,p2425);
HA ha651(p2302,p2304,p2426,p2427);
HA ha652(p2407,p2409,p2428,p2429);
HA ha653(p2411,p2417,p2430,p2431);
FA fa562(p2419,p2423,p2290,p2432,p2433);
HA ha654(p2292,p2306,p2434,p2435);
FA fa563(p2421,p2427,p2429,p2436,p2437);
HA ha655(p2431,p2298,p2438,p2439);
HA ha656(p2300,p2314,p2440,p2441);
FA fa564(p2425,p2433,p2435,p2442,p2443);
FA fa565(p2308,p2310,p2437,p2444,p2445);
HA ha657(p2439,p2441,p2446,p2447);
HA ha658(p2312,p2316,p2448,p2449);
FA fa566(p2443,p2447,p2318,p2450,p2451);
HA ha659(p2445,p2449,p2452,p2453);
FA fa567(p2320,p2322,p2330,p2454,p2455);
HA ha660(p2451,p2453,p2456,p2457);
HA ha661(p2324,p2326,p2458,p2459);
HA ha662(p2328,p2457,p2460,p2461);
HA ha663(p2336,p2455,p2462,p2463);
FA fa568(p2459,p2461,p2332,p2464,p2465);
HA ha664(p2334,p2463,p2466,p2467);
FA fa569(p2465,p2467,p2338,p2468,p2469);
HA ha665(p2340,p2344,p2470,p2471);
HA ha666(p2342,p2346,p2472,p2473);
FA fa570(p2469,p2471,p2473,p2474,p2475);
FA fa571(p2475,p2348,p2350,p2476,p2477);
FA fa572(p2352,p2477,p2354,p2478,p2479);
FA fa573(ip_7_31,ip_8_30,ip_9_29,p2480,p2481);
FA fa574(ip_10_28,ip_11_27,ip_12_26,p2482,p2483);
FA fa575(ip_13_25,ip_14_24,ip_15_23,p2484,p2485);
FA fa576(ip_16_22,ip_17_21,ip_18_20,p2486,p2487);
FA fa577(ip_19_19,ip_20_18,ip_21_17,p2488,p2489);
HA ha667(ip_22_16,ip_23_15,p2490,p2491);
HA ha668(ip_24_14,ip_25_13,p2492,p2493);
HA ha669(ip_26_12,ip_27_11,p2494,p2495);
FA fa578(ip_28_10,ip_29_9,ip_30_8,p2496,p2497);
FA fa579(ip_31_7,p2358,p2360,p2498,p2499);
FA fa580(p2362,p2364,p2366,p2500,p2501);
HA ha670(p2368,p2370,p2502,p2503);
HA ha671(p2372,p2374,p2504,p2505);
HA ha672(p2376,p2378,p2506,p2507);
HA ha673(p2380,p2491,p2508,p2509);
FA fa581(p2493,p2495,p2384,p2510,p2511);
FA fa582(p2386,p2388,p2390,p2512,p2513);
FA fa583(p2392,p2481,p2483,p2514,p2515);
HA ha674(p2485,p2487,p2516,p2517);
HA ha675(p2489,p2497,p2518,p2519);
FA fa584(p2503,p2505,p2507,p2520,p2521);
FA fa585(p2509,p2382,p2400,p2522,p2523);
FA fa586(p2499,p2501,p2511,p2524,p2525);
FA fa587(p2517,p2519,p2394,p2526,p2527);
FA fa588(p2396,p2412,p2414,p2528,p2529);
HA ha676(p2513,p2515,p2530,p2531);
FA fa589(p2521,p2398,p2402,p2532,p2533);
FA fa590(p2404,p2416,p2418,p2534,p2535);
FA fa591(p2422,p2523,p2525,p2536,p2537);
HA ha677(p2527,p2531,p2538,p2539);
FA fa592(p2406,p2408,p2410,p2540,p2541);
FA fa593(p2426,p2428,p2430,p2542,p2543);
HA ha678(p2529,p2539,p2544,p2545);
HA ha679(p2420,p2434,p2546,p2547);
FA fa594(p2533,p2535,p2537,p2548,p2549);
FA fa595(p2545,p2424,p2432,p2550,p2551);
FA fa596(p2438,p2440,p2541,p2552,p2553);
HA ha680(p2543,p2547,p2554,p2555);
FA fa597(p2436,p2446,p2549,p2556,p2557);
FA fa598(p2555,p2442,p2448,p2558,p2559);
FA fa599(p2551,p2553,p2444,p2560,p2561);
FA fa600(p2452,p2557,p2450,p2562,p2563);
HA ha681(p2456,p2559,p2564,p2565);
FA fa601(p2561,p2458,p2460,p2566,p2567);
HA ha682(p2563,p2565,p2568,p2569);
FA fa602(p2454,p2462,p2569,p2570,p2571);
HA ha683(p2466,p2567,p2572,p2573);
FA fa603(p2464,p2571,p2573,p2574,p2575);
HA ha684(p2470,p2468,p2576,p2577);
FA fa604(p2472,p2575,p2577,p2578,p2579);
HA ha685(p2474,p2579,p2580,p2581);
HA ha686(p2581,p2476,p2582,p2583);
HA ha687(ip_8_31,ip_9_30,p2584,p2585);
HA ha688(ip_10_29,ip_11_28,p2586,p2587);
HA ha689(ip_12_27,ip_13_26,p2588,p2589);
HA ha690(ip_14_25,ip_15_24,p2590,p2591);
FA fa605(ip_16_23,ip_17_22,ip_18_21,p2592,p2593);
FA fa606(ip_19_20,ip_20_19,ip_21_18,p2594,p2595);
HA ha691(ip_22_17,ip_23_16,p2596,p2597);
HA ha692(ip_24_15,ip_25_14,p2598,p2599);
HA ha693(ip_26_13,ip_27_12,p2600,p2601);
FA fa607(ip_28_11,ip_29_10,ip_30_9,p2602,p2603);
FA fa608(ip_31_8,p2490,p2492,p2604,p2605);
HA ha694(p2494,p2585,p2606,p2607);
FA fa609(p2587,p2589,p2591,p2608,p2609);
FA fa610(p2597,p2599,p2601,p2610,p2611);
HA ha695(p2502,p2504,p2612,p2613);
FA fa611(p2506,p2508,p2593,p2614,p2615);
HA ha696(p2595,p2603,p2616,p2617);
HA ha697(p2607,p2480,p2618,p2619);
HA ha698(p2482,p2484,p2620,p2621);
FA fa612(p2486,p2488,p2496,p2622,p2623);
FA fa613(p2516,p2518,p2605,p2624,p2625);
FA fa614(p2609,p2611,p2613,p2626,p2627);
HA ha699(p2617,p2498,p2628,p2629);
HA ha700(p2500,p2510,p2630,p2631);
HA ha701(p2615,p2619,p2632,p2633);
FA fa615(p2621,p2512,p2514,p2634,p2635);
FA fa616(p2520,p2530,p2623,p2636,p2637);
FA fa617(p2625,p2627,p2629,p2638,p2639);
FA fa618(p2631,p2633,p2522,p2640,p2641);
HA ha702(p2524,p2526,p2642,p2643);
FA fa619(p2538,p2528,p2544,p2644,p2645);
HA ha703(p2635,p2637,p2646,p2647);
FA fa620(p2639,p2641,p2643,p2648,p2649);
HA ha704(p2532,p2534,p2650,p2651);
FA fa621(p2536,p2546,p2647,p2652,p2653);
FA fa622(p2540,p2542,p2554,p2654,p2655);
HA ha705(p2645,p2649,p2656,p2657);
FA fa623(p2651,p2548,p2653,p2658,p2659);
HA ha706(p2657,p2550,p2660,p2661);
HA ha707(p2552,p2655,p2662,p2663);
FA fa624(p2556,p2659,p2661,p2664,p2665);
FA fa625(p2663,p2558,p2560,p2666,p2667);
FA fa626(p2564,p2562,p2568,p2668,p2669);
HA ha708(p2665,p2667,p2670,p2671);
FA fa627(p2566,p2572,p2669,p2672,p2673);
FA fa628(p2671,p2570,p2673,p2674,p2675);
HA ha709(p2574,p2576,p2676,p2677);
HA ha710(p2675,p2677,p2678,p2679);
HA ha711(p2578,p2580,p2680,p2681);
HA ha712(p2679,p2681,p2682,p2683);
HA ha713(ip_9_31,ip_10_30,p2684,p2685);
HA ha714(ip_11_29,ip_12_28,p2686,p2687);
HA ha715(ip_13_27,ip_14_26,p2688,p2689);
FA fa629(ip_15_25,ip_16_24,ip_17_23,p2690,p2691);
FA fa630(ip_18_22,ip_19_21,ip_20_20,p2692,p2693);
FA fa631(ip_21_19,ip_22_18,ip_23_17,p2694,p2695);
FA fa632(ip_24_16,ip_25_15,ip_26_14,p2696,p2697);
FA fa633(ip_27_13,ip_28_12,ip_29_11,p2698,p2699);
FA fa634(ip_30_10,ip_31_9,p2584,p2700,p2701);
HA ha716(p2586,p2588,p2702,p2703);
FA fa635(p2590,p2596,p2598,p2704,p2705);
HA ha717(p2600,p2685,p2706,p2707);
FA fa636(p2687,p2689,p2606,p2708,p2709);
HA ha718(p2691,p2693,p2710,p2711);
HA ha719(p2695,p2697,p2712,p2713);
FA fa637(p2699,p2701,p2703,p2714,p2715);
HA ha720(p2707,p2592,p2716,p2717);
HA ha721(p2594,p2602,p2718,p2719);
HA ha722(p2612,p2616,p2720,p2721);
HA ha723(p2705,p2709,p2722,p2723);
HA ha724(p2711,p2713,p2724,p2725);
HA ha725(p2604,p2608,p2726,p2727);
HA ha726(p2610,p2618,p2728,p2729);
HA ha727(p2620,p2715,p2730,p2731);
FA fa638(p2717,p2719,p2721,p2732,p2733);
FA fa639(p2723,p2725,p2614,p2734,p2735);
FA fa640(p2628,p2630,p2632,p2736,p2737);
FA fa641(p2727,p2729,p2731,p2738,p2739);
HA ha728(p2622,p2624,p2740,p2741);
FA fa642(p2626,p2733,p2735,p2742,p2743);
FA fa643(p2642,p2737,p2739,p2744,p2745);
FA fa644(p2741,p2634,p2636,p2746,p2747);
HA ha729(p2638,p2640,p2748,p2749);
FA fa645(p2646,p2743,p2650,p2750,p2751);
HA ha730(p2745,p2749,p2752,p2753);
FA fa646(p2644,p2648,p2656,p2754,p2755);
HA ha731(p2747,p2751,p2756,p2757);
HA ha732(p2753,p2652,p2758,p2759);
HA ha733(p2757,p2654,p2760,p2761);
FA fa647(p2660,p2662,p2755,p2762,p2763);
FA fa648(p2759,p2658,p2761,p2764,p2765);
FA fa649(p2763,p2664,p2765,p2766,p2767);
HA ha734(p2666,p2670,p2768,p2769);
FA fa650(p2668,p2767,p2769,p2770,p2771);
HA ha735(p2672,p2771,p2772,p2773);
FA fa651(p2674,p2676,p2773,p2774,p2775);
FA fa652(p2678,p2680,p2775,p2776,p2777);
HA ha736(ip_10_31,ip_11_30,p2778,p2779);
HA ha737(ip_12_29,ip_13_28,p2780,p2781);
FA fa653(ip_14_27,ip_15_26,ip_16_25,p2782,p2783);
HA ha738(ip_17_24,ip_18_23,p2784,p2785);
HA ha739(ip_19_22,ip_20_21,p2786,p2787);
HA ha740(ip_21_20,ip_22_19,p2788,p2789);
HA ha741(ip_23_18,ip_24_17,p2790,p2791);
FA fa654(ip_25_16,ip_26_15,ip_27_14,p2792,p2793);
HA ha742(ip_28_13,ip_29_12,p2794,p2795);
HA ha743(ip_30_11,ip_31_10,p2796,p2797);
FA fa655(p2684,p2686,p2688,p2798,p2799);
HA ha744(p2779,p2781,p2800,p2801);
HA ha745(p2785,p2787,p2802,p2803);
FA fa656(p2789,p2791,p2795,p2804,p2805);
HA ha746(p2797,p2702,p2806,p2807);
HA ha747(p2706,p2783,p2808,p2809);
HA ha748(p2793,p2801,p2810,p2811);
HA ha749(p2803,p2690,p2812,p2813);
HA ha750(p2692,p2694,p2814,p2815);
HA ha751(p2696,p2698,p2816,p2817);
FA fa657(p2700,p2710,p2712,p2818,p2819);
FA fa658(p2799,p2805,p2807,p2820,p2821);
FA fa659(p2809,p2811,p2704,p2822,p2823);
HA ha752(p2708,p2716,p2824,p2825);
HA ha753(p2718,p2720,p2826,p2827);
HA ha754(p2722,p2724,p2828,p2829);
FA fa660(p2813,p2815,p2817,p2830,p2831);
FA fa661(p2714,p2726,p2728,p2832,p2833);
HA ha755(p2730,p2819,p2834,p2835);
HA ha756(p2821,p2823,p2836,p2837);
HA ha757(p2825,p2827,p2838,p2839);
FA fa662(p2829,p2831,p2835,p2840,p2841);
HA ha758(p2837,p2839,p2842,p2843);
FA fa663(p2732,p2734,p2740,p2844,p2845);
FA fa664(p2833,p2843,p2736,p2846,p2847);
HA ha759(p2738,p2841,p2848,p2849);
FA fa665(p2742,p2748,p2845,p2850,p2851);
HA ha760(p2847,p2849,p2852,p2853);
HA ha761(p2744,p2752,p2854,p2855);
HA ha762(p2853,p2746,p2856,p2857);
FA fa666(p2750,p2756,p2851,p2858,p2859);
HA ha763(p2855,p2758,p2860,p2861);
FA fa667(p2857,p2754,p2760,p2862,p2863);
HA ha764(p2859,p2861,p2864,p2865);
FA fa668(p2865,p2762,p2863,p2866,p2867);
HA ha765(p2764,p2768,p2868,p2869);
FA fa669(p2867,p2766,p2869,p2870,p2871);
HA ha766(p2770,p2772,p2872,p2873);
HA ha767(p2871,p2873,p2874,p2875);
HA ha768(p2875,p2774,p2876,p2877);
HA ha769(ip_11_31,ip_12_30,p2878,p2879);
HA ha770(ip_13_29,ip_14_28,p2880,p2881);
HA ha771(ip_15_27,ip_16_26,p2882,p2883);
HA ha772(ip_17_25,ip_18_24,p2884,p2885);
HA ha773(ip_19_23,ip_20_22,p2886,p2887);
FA fa670(ip_21_21,ip_22_20,ip_23_19,p2888,p2889);
FA fa671(ip_24_18,ip_25_17,ip_26_16,p2890,p2891);
HA ha774(ip_27_15,ip_28_14,p2892,p2893);
FA fa672(ip_29_13,ip_30_12,ip_31_11,p2894,p2895);
FA fa673(p2778,p2780,p2784,p2896,p2897);
HA ha775(p2786,p2788,p2898,p2899);
HA ha776(p2790,p2794,p2900,p2901);
HA ha777(p2796,p2879,p2902,p2903);
HA ha778(p2881,p2883,p2904,p2905);
HA ha779(p2885,p2887,p2906,p2907);
FA fa674(p2893,p2800,p2802,p2908,p2909);
FA fa675(p2889,p2891,p2895,p2910,p2911);
HA ha780(p2899,p2901,p2912,p2913);
HA ha781(p2903,p2905,p2914,p2915);
FA fa676(p2907,p2782,p2792,p2916,p2917);
FA fa677(p2806,p2808,p2810,p2918,p2919);
HA ha782(p2897,p2913,p2920,p2921);
HA ha783(p2915,p2798,p2922,p2923);
HA ha784(p2804,p2812,p2924,p2925);
HA ha785(p2814,p2816,p2926,p2927);
FA fa678(p2909,p2911,p2921,p2928,p2929);
FA fa679(p2824,p2826,p2828,p2930,p2931);
HA ha786(p2917,p2919,p2932,p2933);
FA fa680(p2923,p2925,p2927,p2934,p2935);
HA ha787(p2818,p2820,p2936,p2937);
FA fa681(p2822,p2834,p2836,p2938,p2939);
FA fa682(p2838,p2929,p2933,p2940,p2941);
FA fa683(p2830,p2842,p2931,p2942,p2943);
HA ha788(p2935,p2937,p2944,p2945);
FA fa684(p2832,p2939,p2941,p2946,p2947);
FA fa685(p2945,p2840,p2848,p2948,p2949);
HA ha789(p2943,p2844,p2950,p2951);
FA fa686(p2846,p2852,p2947,p2952,p2953);
FA fa687(p2854,p2949,p2951,p2954,p2955);
HA ha790(p2850,p2856,p2956,p2957);
FA fa688(p2953,p2860,p2955,p2958,p2959);
FA fa689(p2957,p2858,p2864,p2960,p2961);
HA ha791(p2959,p2862,p2962,p2963);
HA ha792(p2961,p2963,p2964,p2965);
HA ha793(p2866,p2868,p2966,p2967);
HA ha794(p2965,p2967,p2968,p2969);
HA ha795(p2969,p2870,p2970,p2971);
HA ha796(p2872,p2874,p2972,p2973);
HA ha797(p2971,p2973,p2974,p2975);
HA ha798(ip_12_31,ip_13_30,p2976,p2977);
HA ha799(ip_14_29,ip_15_28,p2978,p2979);
HA ha800(ip_16_27,ip_17_26,p2980,p2981);
FA fa690(ip_18_25,ip_19_24,ip_20_23,p2982,p2983);
HA ha801(ip_21_22,ip_22_21,p2984,p2985);
FA fa691(ip_23_20,ip_24_19,ip_25_18,p2986,p2987);
FA fa692(ip_26_17,ip_27_16,ip_28_15,p2988,p2989);
FA fa693(ip_29_14,ip_30_13,ip_31_12,p2990,p2991);
HA ha802(p2878,p2880,p2992,p2993);
FA fa694(p2882,p2884,p2886,p2994,p2995);
HA ha803(p2892,p2977,p2996,p2997);
HA ha804(p2979,p2981,p2998,p2999);
FA fa695(p2985,p2898,p2900,p3000,p3001);
HA ha805(p2902,p2904,p3002,p3003);
HA ha806(p2906,p2983,p3004,p3005);
FA fa696(p2987,p2989,p2991,p3006,p3007);
HA ha807(p2993,p2997,p3008,p3009);
HA ha808(p2999,p2888,p3010,p3011);
FA fa697(p2890,p2894,p2912,p3012,p3013);
HA ha809(p2914,p2995,p3014,p3015);
HA ha810(p3003,p3005,p3016,p3017);
FA fa698(p3009,p2896,p2920,p3018,p3019);
FA fa699(p3001,p3007,p3011,p3020,p3021);
HA ha811(p3015,p3017,p3022,p3023);
FA fa700(p2908,p2910,p2922,p3024,p3025);
FA fa701(p2924,p2926,p3013,p3026,p3027);
FA fa702(p3023,p2916,p2918,p3028,p3029);
FA fa703(p2932,p3019,p3021,p3030,p3031);
FA fa704(p2928,p2936,p3025,p3032,p3033);
HA ha812(p3027,p2930,p3034,p3035);
HA ha813(p2934,p2944,p3036,p3037);
HA ha814(p3029,p3031,p3038,p3039);
HA ha815(p2938,p2940,p3040,p3041);
HA ha816(p3033,p3035,p3042,p3043);
HA ha817(p3037,p3039,p3044,p3045);
FA fa705(p2942,p3041,p3043,p3046,p3047);
FA fa706(p3045,p2946,p2950,p3048,p3049);
FA fa707(p2948,p3047,p2952,p3050,p3051);
HA ha818(p2956,p3049,p3052,p3053);
FA fa708(p2954,p3051,p3053,p3054,p3055);
FA fa709(p2958,p3055,p2960,p3056,p3057);
HA ha819(p2962,p2964,p3058,p3059);
FA fa710(p3057,p2966,p3059,p3060,p3061);
FA fa711(p2968,p3061,p2970,p3062,p3063);
FA fa712(p2972,p3063,p2974,p3064,p3065);
HA ha820(ip_13_31,ip_14_30,p3066,p3067);
FA fa713(ip_15_29,ip_16_28,ip_17_27,p3068,p3069);
HA ha821(ip_18_26,ip_19_25,p3070,p3071);
HA ha822(ip_20_24,ip_21_23,p3072,p3073);
FA fa714(ip_22_22,ip_23_21,ip_24_20,p3074,p3075);
HA ha823(ip_25_19,ip_26_18,p3076,p3077);
HA ha824(ip_27_17,ip_28_16,p3078,p3079);
FA fa715(ip_29_15,ip_30_14,ip_31_13,p3080,p3081);
FA fa716(p2976,p2978,p2980,p3082,p3083);
FA fa717(p2984,p3067,p3071,p3084,p3085);
FA fa718(p3073,p3077,p3079,p3086,p3087);
FA fa719(p2992,p2996,p2998,p3088,p3089);
HA ha825(p3069,p3075,p3090,p3091);
HA ha826(p3081,p2982,p3092,p3093);
HA ha827(p2986,p2988,p3094,p3095);
FA fa720(p2990,p3002,p3004,p3096,p3097);
HA ha828(p3008,p3083,p3098,p3099);
HA ha829(p3085,p3087,p3100,p3101);
FA fa721(p3091,p2994,p3010,p3102,p3103);
HA ha830(p3014,p3016,p3104,p3105);
HA ha831(p3089,p3093,p3106,p3107);
HA ha832(p3095,p3099,p3108,p3109);
FA fa722(p3101,p3000,p3006,p3110,p3111);
HA ha833(p3022,p3097,p3112,p3113);
HA ha834(p3105,p3107,p3114,p3115);
FA fa723(p3109,p3012,p3103,p3116,p3117);
HA ha835(p3113,p3115,p3118,p3119);
FA fa724(p3018,p3020,p3111,p3120,p3121);
HA ha836(p3119,p3024,p3122,p3123);
FA fa725(p3026,p3117,p3028,p3124,p3125);
FA fa726(p3030,p3034,p3036,p3126,p3127);
HA ha837(p3038,p3121,p3128,p3129);
HA ha838(p3123,p3032,p3130,p3131);
HA ha839(p3040,p3042,p3132,p3133);
FA fa727(p3044,p3125,p3129,p3134,p3135);
HA ha840(p3127,p3131,p3136,p3137);
HA ha841(p3133,p3135,p3138,p3139);
FA fa728(p3137,p3046,p3139,p3140,p3141);
HA ha842(p3048,p3052,p3142,p3143);
HA ha843(p3050,p3141,p3144,p3145);
HA ha844(p3143,p3145,p3146,p3147);
FA fa729(p3054,p3147,p3056,p3148,p3149);
FA fa730(p3058,p3149,p3060,p3150,p3151);
HA ha845(p3151,p3062,p3152,p3153);
HA ha846(ip_14_31,ip_15_30,p3154,p3155);
FA fa731(ip_16_29,ip_17_28,ip_18_27,p3156,p3157);
FA fa732(ip_19_26,ip_20_25,ip_21_24,p3158,p3159);
HA ha847(ip_22_23,ip_23_22,p3160,p3161);
FA fa733(ip_24_21,ip_25_20,ip_26_19,p3162,p3163);
FA fa734(ip_27_18,ip_28_17,ip_29_16,p3164,p3165);
HA ha848(ip_30_15,ip_31_14,p3166,p3167);
HA ha849(p3066,p3070,p3168,p3169);
FA fa735(p3072,p3076,p3078,p3170,p3171);
HA ha850(p3155,p3161,p3172,p3173);
HA ha851(p3167,p3157,p3174,p3175);
HA ha852(p3159,p3163,p3176,p3177);
HA ha853(p3165,p3169,p3178,p3179);
HA ha854(p3173,p3068,p3180,p3181);
HA ha855(p3074,p3080,p3182,p3183);
HA ha856(p3090,p3171,p3184,p3185);
HA ha857(p3175,p3177,p3186,p3187);
FA fa736(p3179,p3082,p3084,p3188,p3189);
FA fa737(p3086,p3092,p3094,p3190,p3191);
FA fa738(p3098,p3100,p3181,p3192,p3193);
HA ha858(p3183,p3185,p3194,p3195);
FA fa739(p3187,p3088,p3104,p3196,p3197);
HA ha859(p3106,p3108,p3198,p3199);
HA ha860(p3195,p3096,p3200,p3201);
FA fa740(p3112,p3114,p3189,p3202,p3203);
FA fa741(p3191,p3193,p3199,p3204,p3205);
HA ha861(p3102,p3118,p3206,p3207);
FA fa742(p3197,p3201,p3110,p3208,p3209);
FA fa743(p3203,p3205,p3207,p3210,p3211);
HA ha862(p3116,p3122,p3212,p3213);
FA fa744(p3209,p3120,p3128,p3214,p3215);
HA ha863(p3211,p3213,p3216,p3217);
HA ha864(p3124,p3130,p3218,p3219);
HA ha865(p3132,p3217,p3220,p3221);
FA fa745(p3126,p3136,p3215,p3222,p3223);
HA ha866(p3219,p3221,p3224,p3225);
HA ha867(p3134,p3138,p3226,p3227);
FA fa746(p3225,p3223,p3227,p3228,p3229);
FA fa747(p3142,p3140,p3144,p3230,p3231);
FA fa748(p3229,p3146,p3231,p3232,p3233);
FA fa749(p3233,p3148,p3150,p3234,p3235);
HA ha868(ip_15_31,ip_16_30,p3236,p3237);
FA fa750(ip_17_29,ip_18_28,ip_19_27,p3238,p3239);
FA fa751(ip_20_26,ip_21_25,ip_22_24,p3240,p3241);
FA fa752(ip_23_23,ip_24_22,ip_25_21,p3242,p3243);
FA fa753(ip_26_20,ip_27_19,ip_28_18,p3244,p3245);
HA ha869(ip_29_17,ip_30_16,p3246,p3247);
HA ha870(ip_31_15,p3154,p3248,p3249);
FA fa754(p3160,p3166,p3237,p3250,p3251);
FA fa755(p3247,p3168,p3172,p3252,p3253);
HA ha871(p3239,p3241,p3254,p3255);
HA ha872(p3243,p3245,p3256,p3257);
FA fa756(p3249,p3156,p3158,p3258,p3259);
FA fa757(p3162,p3164,p3174,p3260,p3261);
HA ha873(p3176,p3178,p3262,p3263);
HA ha874(p3251,p3255,p3264,p3265);
FA fa758(p3257,p3170,p3180,p3266,p3267);
HA ha875(p3182,p3184,p3268,p3269);
HA ha876(p3186,p3253,p3270,p3271);
FA fa759(p3263,p3265,p3194,p3272,p3273);
HA ha877(p3259,p3261,p3274,p3275);
FA fa760(p3269,p3271,p3198,p3276,p3277);
HA ha878(p3267,p3273,p3278,p3279);
HA ha879(p3275,p3188,p3280,p3281);
HA ha880(p3190,p3192,p3282,p3283);
HA ha881(p3200,p3277,p3284,p3285);
HA ha882(p3279,p3196,p3286,p3287);
HA ha883(p3206,p3281,p3288,p3289);
HA ha884(p3283,p3285,p3290,p3291);
FA fa761(p3202,p3204,p3287,p3292,p3293);
HA ha885(p3289,p3291,p3294,p3295);
HA ha886(p3208,p3212,p3296,p3297);
HA ha887(p3295,p3210,p3298,p3299);
FA fa762(p3216,p3293,p3297,p3300,p3301);
FA fa763(p3218,p3220,p3299,p3302,p3303);
HA ha888(p3214,p3224,p3304,p3305);
HA ha889(p3301,p3226,p3306,p3307);
HA ha890(p3303,p3305,p3308,p3309);
FA fa764(p3222,p3307,p3309,p3310,p3311);
FA fa765(p3228,p3311,p3230,p3312,p3313);
FA fa766(p3232,p3313,p3234,p3314,p3315);
FA fa767(ip_16_31,ip_17_30,ip_18_29,p3316,p3317);
HA ha891(ip_19_28,ip_20_27,p3318,p3319);
FA fa768(ip_21_26,ip_22_25,ip_23_24,p3320,p3321);
FA fa769(ip_24_23,ip_25_22,ip_26_21,p3322,p3323);
HA ha892(ip_27_20,ip_28_19,p3324,p3325);
FA fa770(ip_29_18,ip_30_17,ip_31_16,p3326,p3327);
HA ha893(p3236,p3246,p3328,p3329);
FA fa771(p3319,p3325,p3248,p3330,p3331);
FA fa772(p3317,p3321,p3323,p3332,p3333);
HA ha894(p3327,p3329,p3334,p3335);
HA ha895(p3238,p3240,p3336,p3337);
HA ha896(p3242,p3244,p3338,p3339);
FA fa773(p3254,p3256,p3331,p3340,p3341);
FA fa774(p3335,p3250,p3262,p3342,p3343);
FA fa775(p3264,p3333,p3337,p3344,p3345);
FA fa776(p3339,p3252,p3268,p3346,p3347);
FA fa777(p3270,p3341,p3258,p3348,p3349);
FA fa778(p3260,p3274,p3343,p3350,p3351);
HA ha897(p3345,p3266,p3352,p3353);
FA fa779(p3272,p3278,p3347,p3354,p3355);
FA fa780(p3349,p3276,p3280,p3356,p3357);
HA ha898(p3282,p3284,p3358,p3359);
HA ha899(p3351,p3353,p3360,p3361);
HA ha900(p3286,p3288,p3362,p3363);
HA ha901(p3290,p3355,p3364,p3365);
FA fa781(p3359,p3361,p3294,p3366,p3367);
FA fa782(p3357,p3363,p3365,p3368,p3369);
FA fa783(p3296,p3367,p3292,p3370,p3371);
HA ha902(p3298,p3369,p3372,p3373);
HA ha903(p3371,p3373,p3374,p3375);
FA fa784(p3300,p3304,p3375,p3376,p3377);
HA ha904(p3302,p3306,p3378,p3379);
FA fa785(p3308,p3377,p3379,p3380,p3381);
FA fa786(p3310,p3381,p3312,p3382,p3383);
HA ha905(ip_17_31,ip_18_30,p3384,p3385);
HA ha906(ip_19_29,ip_20_28,p3386,p3387);
HA ha907(ip_21_27,ip_22_26,p3388,p3389);
HA ha908(ip_23_25,ip_24_24,p3390,p3391);
HA ha909(ip_25_23,ip_26_22,p3392,p3393);
FA fa787(ip_27_21,ip_28_20,ip_29_19,p3394,p3395);
HA ha910(ip_30_18,ip_31_17,p3396,p3397);
HA ha911(p3318,p3324,p3398,p3399);
FA fa788(p3385,p3387,p3389,p3400,p3401);
FA fa789(p3391,p3393,p3397,p3402,p3403);
HA ha912(p3328,p3395,p3404,p3405);
FA fa790(p3399,p3316,p3320,p3406,p3407);
FA fa791(p3322,p3326,p3334,p3408,p3409);
HA ha913(p3401,p3403,p3410,p3411);
HA ha914(p3405,p3330,p3412,p3413);
FA fa792(p3336,p3338,p3411,p3414,p3415);
HA ha915(p3332,p3407,p3416,p3417);
HA ha916(p3409,p3413,p3418,p3419);
FA fa793(p3340,p3415,p3417,p3420,p3421);
HA ha917(p3419,p3342,p3422,p3423);
HA ha918(p3344,p3346,p3424,p3425);
HA ha919(p3348,p3352,p3426,p3427);
HA ha920(p3421,p3423,p3428,p3429);
FA fa794(p3350,p3358,p3360,p3430,p3431);
FA fa795(p3425,p3427,p3429,p3432,p3433);
HA ha921(p3354,p3362,p3434,p3435);
HA ha922(p3364,p3356,p3436,p3437);
HA ha923(p3431,p3433,p3438,p3439);
HA ha924(p3435,p3366,p3440,p3441);
HA ha925(p3437,p3439,p3442,p3443);
FA fa796(p3368,p3372,p3441,p3444,p3445);
HA ha926(p3443,p3370,p3446,p3447);
FA fa797(p3374,p3445,p3447,p3448,p3449);
FA fa798(p3378,p3376,p3449,p3450,p3451);
FA fa799(p3380,p3451,p3382,p3452,p3453);
HA ha927(ip_18_31,ip_19_30,p3454,p3455);
FA fa800(ip_20_29,ip_21_28,ip_22_27,p3456,p3457);
FA fa801(ip_23_26,ip_24_25,ip_25_24,p3458,p3459);
HA ha928(ip_26_23,ip_27_22,p3460,p3461);
FA fa802(ip_28_21,ip_29_20,ip_30_19,p3462,p3463);
FA fa803(ip_31_18,p3384,p3386,p3464,p3465);
HA ha929(p3388,p3390,p3466,p3467);
FA fa804(p3392,p3396,p3455,p3468,p3469);
HA ha930(p3461,p3398,p3470,p3471);
HA ha931(p3457,p3459,p3472,p3473);
FA fa805(p3463,p3467,p3394,p3474,p3475);
HA ha932(p3404,p3465,p3476,p3477);
FA fa806(p3469,p3471,p3473,p3478,p3479);
FA fa807(p3400,p3402,p3410,p3480,p3481);
FA fa808(p3475,p3477,p3412,p3482,p3483);
HA ha933(p3479,p3406,p3484,p3485);
FA fa809(p3408,p3416,p3418,p3486,p3487);
FA fa810(p3481,p3483,p3414,p3488,p3489);
HA ha934(p3485,p3422,p3490,p3491);
HA ha935(p3487,p3489,p3492,p3493);
FA fa811(p3420,p3424,p3426,p3494,p3495);
HA ha936(p3428,p3491,p3496,p3497);
FA fa812(p3493,p3497,p3434,p3498,p3499);
FA fa813(p3495,p3430,p3432,p3500,p3501);
FA fa814(p3436,p3438,p3499,p3502,p3503);
FA fa815(p3440,p3442,p3501,p3504,p3505);
FA fa816(p3503,p3446,p3505,p3506,p3507);
HA ha937(p3444,p3507,p3508,p3509);
HA ha938(p3448,p3509,p3510,p3511);
FA fa817(p3511,p3450,p3452,p3512,p3513);
FA fa818(ip_19_31,ip_20_30,ip_21_29,p3514,p3515);
HA ha939(ip_22_28,ip_23_27,p3516,p3517);
HA ha940(ip_24_26,ip_25_25,p3518,p3519);
FA fa819(ip_26_24,ip_27_23,ip_28_22,p3520,p3521);
FA fa820(ip_29_21,ip_30_20,ip_31_19,p3522,p3523);
HA ha941(p3454,p3460,p3524,p3525);
HA ha942(p3517,p3519,p3526,p3527);
FA fa821(p3466,p3515,p3521,p3528,p3529);
HA ha943(p3523,p3525,p3530,p3531);
HA ha944(p3527,p3456,p3532,p3533);
FA fa822(p3458,p3462,p3470,p3534,p3535);
HA ha945(p3472,p3531,p3536,p3537);
FA fa823(p3464,p3468,p3476,p3538,p3539);
FA fa824(p3529,p3533,p3537,p3540,p3541);
HA ha946(p3474,p3535,p3542,p3543);
FA fa825(p3478,p3539,p3541,p3544,p3545);
HA ha947(p3543,p3480,p3546,p3547);
HA ha948(p3482,p3484,p3548,p3549);
FA fa826(p3545,p3547,p3549,p3550,p3551);
FA fa827(p3486,p3488,p3490,p3552,p3553);
HA ha949(p3492,p3496,p3554,p3555);
HA ha950(p3551,p3553,p3556,p3557);
HA ha951(p3555,p3494,p3558,p3559);
HA ha952(p3557,p3498,p3560,p3561);
HA ha953(p3559,p3561,p3562,p3563);
HA ha954(p3500,p3502,p3564,p3565);
FA fa828(p3563,p3504,p3565,p3566,p3567);
HA ha955(p3506,p3508,p3568,p3569);
FA fa829(p3567,p3510,p3569,p3570,p3571);
HA ha956(ip_20_31,ip_21_30,p3572,p3573);
HA ha957(ip_22_29,ip_23_28,p3574,p3575);
FA fa830(ip_24_27,ip_25_26,ip_26_25,p3576,p3577);
FA fa831(ip_27_24,ip_28_23,ip_29_22,p3578,p3579);
FA fa832(ip_30_21,ip_31_20,p3516,p3580,p3581);
FA fa833(p3518,p3573,p3575,p3582,p3583);
HA ha958(p3524,p3526,p3584,p3585);
HA ha959(p3577,p3579,p3586,p3587);
FA fa834(p3581,p3514,p3520,p3588,p3589);
FA fa835(p3522,p3530,p3583,p3590,p3591);
HA ha960(p3585,p3587,p3592,p3593);
HA ha961(p3532,p3536,p3594,p3595);
HA ha962(p3593,p3528,p3596,p3597);
HA ha963(p3589,p3591,p3598,p3599);
HA ha964(p3595,p3534,p3600,p3601);
FA fa836(p3542,p3597,p3599,p3602,p3603);
FA fa837(p3538,p3540,p3601,p3604,p3605);
HA ha965(p3546,p3548,p3606,p3607);
FA fa838(p3603,p3544,p3605,p3608,p3609);
FA fa839(p3607,p3550,p3554,p3610,p3611);
HA ha966(p3609,p3552,p3612,p3613);
HA ha967(p3556,p3558,p3614,p3615);
FA fa840(p3611,p3613,p3560,p3616,p3617);
FA fa841(p3615,p3562,p3617,p3618,p3619);
HA ha968(p3564,p3619,p3620,p3621);
HA ha969(p3621,p3566,p3622,p3623);
HA ha970(p3568,p3623,p3624,p3625);
FA fa842(ip_21_31,ip_22_30,ip_23_29,p3626,p3627);
HA ha971(ip_24_28,ip_25_27,p3628,p3629);
HA ha972(ip_26_26,ip_27_25,p3630,p3631);
HA ha973(ip_28_24,ip_29_23,p3632,p3633);
HA ha974(ip_30_22,ip_31_21,p3634,p3635);
FA fa843(p3572,p3574,p3629,p3636,p3637);
FA fa844(p3631,p3633,p3635,p3638,p3639);
FA fa845(p3627,p3576,p3578,p3640,p3641);
HA ha975(p3580,p3584,p3642,p3643);
FA fa846(p3586,p3637,p3639,p3644,p3645);
HA ha976(p3582,p3592,p3646,p3647);
HA ha977(p3643,p3594,p3648,p3649);
FA fa847(p3641,p3645,p3647,p3650,p3651);
FA fa848(p3588,p3590,p3596,p3652,p3653);
HA ha978(p3598,p3649,p3654,p3655);
FA fa849(p3600,p3651,p3655,p3656,p3657);
FA fa850(p3653,p3602,p3606,p3658,p3659);
HA ha979(p3657,p3604,p3660,p3661);
HA ha980(p3659,p3661,p3662,p3663);
HA ha981(p3608,p3663,p3664,p3665);
FA fa851(p3612,p3665,p3610,p3666,p3667);
HA ha982(p3614,p3667,p3668,p3669);
FA fa852(p3616,p3669,p3618,p3670,p3671);
FA fa853(p3620,p3671,p3622,p3672,p3673);
HA ha983(ip_22_31,ip_23_30,p3674,p3675);
HA ha984(ip_24_29,ip_25_28,p3676,p3677);
HA ha985(ip_26_27,ip_27_26,p3678,p3679);
FA fa854(ip_28_25,ip_29_24,ip_30_23,p3680,p3681);
HA ha986(ip_31_22,p3628,p3682,p3683);
FA fa855(p3630,p3632,p3634,p3684,p3685);
FA fa856(p3675,p3677,p3679,p3686,p3687);
FA fa857(p3681,p3683,p3626,p3688,p3689);
FA fa858(p3685,p3687,p3636,p3690,p3691);
HA ha987(p3638,p3642,p3692,p3693);
FA fa859(p3689,p3646,p3691,p3694,p3695);
FA fa860(p3693,p3640,p3644,p3696,p3697);
FA fa861(p3648,p3654,p3695,p3698,p3699);
HA ha988(p3650,p3697,p3700,p3701);
FA fa862(p3652,p3699,p3701,p3702,p3703);
HA ha989(p3656,p3660,p3704,p3705);
HA ha990(p3703,p3658,p3706,p3707);
FA fa863(p3662,p3705,p3664,p3708,p3709);
HA ha991(p3707,p3709,p3710,p3711);
HA ha992(p3711,p3666,p3712,p3713);
FA fa864(p3668,p3713,p3670,p3714,p3715);
HA ha993(ip_23_31,ip_24_30,p3716,p3717);
HA ha994(ip_25_29,ip_26_28,p3718,p3719);
HA ha995(ip_27_27,ip_28_26,p3720,p3721);
HA ha996(ip_29_25,ip_30_24,p3722,p3723);
HA ha997(ip_31_23,p3674,p3724,p3725);
HA ha998(p3676,p3678,p3726,p3727);
FA fa865(p3717,p3719,p3721,p3728,p3729);
HA ha999(p3723,p3682,p3730,p3731);
HA ha1000(p3725,p3727,p3732,p3733);
HA ha1001(p3680,p3729,p3734,p3735);
HA ha1002(p3731,p3733,p3736,p3737);
FA fa866(p3684,p3686,p3735,p3738,p3739);
HA ha1003(p3737,p3688,p3740,p3741);
HA ha1004(p3692,p3690,p3742,p3743);
FA fa867(p3739,p3741,p3743,p3744,p3745);
FA fa868(p3694,p3745,p3696,p3746,p3747);
HA ha1005(p3700,p3698,p3748,p3749);
FA fa869(p3747,p3749,p3702,p3750,p3751);
FA fa870(p3704,p3706,p3751,p3752,p3753);
HA ha1006(p3708,p3710,p3754,p3755);
HA ha1007(p3753,p3755,p3756,p3757);
HA ha1008(p3712,p3757,p3758,p3759);
HA ha1009(ip_24_31,ip_25_30,p3760,p3761);
HA ha1010(ip_26_29,ip_27_28,p3762,p3763);
HA ha1011(ip_28_27,ip_29_26,p3764,p3765);
HA ha1012(ip_30_25,ip_31_24,p3766,p3767);
HA ha1013(p3716,p3718,p3768,p3769);
HA ha1014(p3720,p3722,p3770,p3771);
HA ha1015(p3761,p3763,p3772,p3773);
HA ha1016(p3765,p3767,p3774,p3775);
HA ha1017(p3724,p3726,p3776,p3777);
HA ha1018(p3769,p3771,p3778,p3779);
FA fa871(p3773,p3775,p3730,p3780,p3781);
FA fa872(p3732,p3777,p3779,p3782,p3783);
HA ha1019(p3728,p3734,p3784,p3785);
HA ha1020(p3736,p3781,p3786,p3787);
FA fa873(p3783,p3785,p3787,p3788,p3789);
HA ha1021(p3740,p3738,p3790,p3791);
HA ha1022(p3742,p3789,p3792,p3793);
HA ha1023(p3791,p3793,p3794,p3795);
HA ha1024(p3744,p3795,p3796,p3797);
HA ha1025(p3797,p3746,p3798,p3799);
HA ha1026(p3748,p3799,p3800,p3801);
FA fa874(p3801,p3750,p3752,p3802,p3803);
FA fa875(p3754,p3756,p3803,p3804,p3805);
HA ha1027(ip_25_31,ip_26_30,p3806,p3807);
HA ha1028(ip_27_29,ip_28_28,p3808,p3809);
HA ha1029(ip_29_27,ip_30_26,p3810,p3811);
HA ha1030(ip_31_25,p3760,p3812,p3813);
FA fa876(p3762,p3764,p3766,p3814,p3815);
FA fa877(p3807,p3809,p3811,p3816,p3817);
FA fa878(p3768,p3770,p3772,p3818,p3819);
HA ha1031(p3774,p3813,p3820,p3821);
FA fa879(p3776,p3778,p3815,p3822,p3823);
HA ha1032(p3817,p3821,p3824,p3825);
HA ha1033(p3819,p3825,p3826,p3827);
HA ha1034(p3780,p3784,p3828,p3829);
HA ha1035(p3786,p3823,p3830,p3831);
FA fa880(p3827,p3782,p3829,p3832,p3833);
FA fa881(p3831,p3788,p3790,p3834,p3835);
HA ha1036(p3792,p3833,p3836,p3837);
HA ha1037(p3794,p3837,p3838,p3839);
HA ha1038(p3796,p3835,p3840,p3841);
HA ha1039(p3839,p3841,p3842,p3843);
HA ha1040(p3798,p3843,p3844,p3845);
FA fa882(p3800,p3845,p3802,p3846,p3847);
HA ha1041(ip_26_31,ip_27_30,p3848,p3849);
FA fa883(ip_28_29,ip_29_28,ip_30_27,p3850,p3851);
HA ha1042(ip_31_26,p3806,p3852,p3853);
HA ha1043(p3808,p3810,p3854,p3855);
HA ha1044(p3849,p3812,p3856,p3857);
HA ha1045(p3851,p3853,p3858,p3859);
FA fa884(p3855,p3820,p3857,p3860,p3861);
HA ha1046(p3859,p3814,p3862,p3863);
FA fa885(p3816,p3824,p3818,p3864,p3865);
HA ha1047(p3826,p3861,p3866,p3867);
FA fa886(p3863,p3822,p3828,p3868,p3869);
HA ha1048(p3830,p3865,p3870,p3871);
HA ha1049(p3867,p3871,p3872,p3873);
FA fa887(p3869,p3873,p3832,p3874,p3875);
HA ha1050(p3836,p3838,p3876,p3877);
HA ha1051(p3875,p3834,p3878,p3879);
FA fa888(p3840,p3877,p3842,p3880,p3881);
HA ha1052(p3879,p3844,p3882,p3883);
FA fa889(p3881,p3883,p3846,p3884,p3885);
HA ha1053(ip_27_31,ip_28_30,p3886,p3887);
HA ha1054(ip_29_29,ip_30_28,p3888,p3889);
HA ha1055(ip_31_27,p3848,p3890,p3891);
FA fa890(p3887,p3889,p3852,p3892,p3893);
HA ha1056(p3854,p3891,p3894,p3895);
HA ha1057(p3850,p3856,p3896,p3897);
HA ha1058(p3858,p3893,p3898,p3899);
HA ha1059(p3895,p3897,p3900,p3901);
HA ha1060(p3899,p3862,p3902,p3903);
FA fa891(p3901,p3860,p3866,p3904,p3905);
FA fa892(p3903,p3864,p3870,p3906,p3907);
HA ha1061(p3872,p3905,p3908,p3909);
FA fa893(p3868,p3907,p3909,p3910,p3911);
FA fa894(p3874,p3876,p3911,p3912,p3913);
HA ha1062(p3878,p3913,p3914,p3915);
FA fa895(p3880,p3882,p3915,p3916,p3917);
HA ha1063(ip_28_31,ip_29_30,p3918,p3919);
FA fa896(ip_30_29,ip_31_28,p3886,p3920,p3921);
HA ha1064(p3888,p3919,p3922,p3923);
FA fa897(p3890,p3921,p3923,p3924,p3925);
FA fa898(p3894,p3892,p3896,p3926,p3927);
FA fa899(p3898,p3925,p3900,p3928,p3929);
HA ha1065(p3902,p3927,p3930,p3931);
HA ha1066(p3929,p3931,p3932,p3933);
HA ha1067(p3933,p3904,p3934,p3935);
FA fa900(p3908,p3906,p3935,p3936,p3937);
FA fa901(p3910,p3937,p3912,p3938,p3939);
HA ha1068(p3914,p3939,p3940,p3941);
FA fa902(ip_29_31,ip_30_30,ip_31_29,p3942,p3943);
HA ha1069(p3918,p3922,p3944,p3945);
FA fa903(p3943,p3920,p3945,p3946,p3947);
HA ha1070(p3924,p3947,p3948,p3949);
HA ha1071(p3949,p3926,p3950,p3951);
HA ha1072(p3928,p3930,p3952,p3953);
HA ha1073(p3932,p3951,p3954,p3955);
FA fa904(p3953,p3955,p3934,p3956,p3957);
FA fa905(p3957,p3936,p3938,p3958,p3959);
HA ha1074(ip_30_31,ip_31_30,p3960,p3961);
FA fa906(p3961,p3942,p3944,p3962,p3963);
FA fa907(p3963,p3946,p3948,p3964,p3965);
HA ha1075(p3950,p3952,p3966,p3967);
FA fa908(p3965,p3954,p3967,p3968,p3969);
FA fa909(p3969,p3956,p3958,p3970,p3971);
FA fa910(ip_31_31,p3960,p3962,p3972,p3973);
FA fa911(p3973,p3964,p3966,p3974,p3975);
HA ha1076(p3975,p3968,p3976,p3977);
wire [63:0] a,b;
wire [63:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p0;
assign b[3] = p5;
assign a[4] = p4;
assign b[4] = p11;
assign a[5] = p19;
assign b[5] = 1'b0;
assign a[6] = p33;
assign b[6] = p18;
assign a[7] = p49;
assign b[7] = p51;
assign a[8] = p50;
assign b[8] = p71;
assign a[9] = p95;
assign b[9] = 1'b0;
assign a[10] = p121;
assign b[10] = p94;
assign a[11] = p120;
assign b[11] = p149;
assign a[12] = p181;
assign b[12] = p148;
assign a[13] = p219;
assign b[13] = p221;
assign a[14] = p265;
assign b[14] = p267;
assign a[15] = p315;
assign b[15] = p317;
assign a[16] = p373;
assign b[16] = 1'b0;
assign a[17] = p429;
assign b[17] = 1'b0;
assign a[18] = p491;
assign b[18] = 1'b0;
assign a[19] = p551;
assign b[19] = p490;
assign a[20] = p619;
assign b[20] = p550;
assign a[21] = p618;
assign b[21] = p687;
assign a[22] = p763;
assign b[22] = 1'b0;
assign a[23] = p849;
assign b[23] = p762;
assign a[24] = p848;
assign b[24] = p933;
assign a[25] = p1025;
assign b[25] = 1'b0;
assign a[26] = p1127;
assign b[26] = p1024;
assign a[27] = p1225;
assign b[27] = p1126;
assign a[28] = p1329;
assign b[28] = p1331;
assign a[29] = p1451;
assign b[29] = p1453;
assign a[30] = p1452;
assign b[30] = p1583;
assign a[31] = p1711;
assign b[31] = 1'b0;
assign a[32] = p1841;
assign b[32] = p1710;
assign a[33] = p1975;
assign b[33] = p1840;
assign a[34] = p2107;
assign b[34] = 1'b0;
assign a[35] = p2239;
assign b[35] = p2106;
assign a[36] = p2238;
assign b[36] = p2357;
assign a[37] = p2479;
assign b[37] = p2356;
assign a[38] = p2583;
assign b[38] = p2478;
assign a[39] = p2683;
assign b[39] = p2582;
assign a[40] = p2682;
assign b[40] = p2777;
assign a[41] = p2877;
assign b[41] = p2776;
assign a[42] = p2876;
assign b[42] = p2975;
assign a[43] = p3065;
assign b[43] = 1'b0;
assign a[44] = p3153;
assign b[44] = p3064;
assign a[45] = p3152;
assign b[45] = p3235;
assign a[46] = p3315;
assign b[46] = 1'b0;
assign a[47] = p3383;
assign b[47] = p3314;
assign a[48] = p3453;
assign b[48] = 1'b0;
assign a[49] = p3513;
assign b[49] = 1'b0;
assign a[50] = p3571;
assign b[50] = p3512;
assign a[51] = p3625;
assign b[51] = p3570;
assign a[52] = p3624;
assign b[52] = p3673;
assign a[53] = p3715;
assign b[53] = p3672;
assign a[54] = p3759;
assign b[54] = p3714;
assign a[55] = p3758;
assign b[55] = p3805;
assign a[56] = p3847;
assign b[56] = p3804;
assign a[57] = p3885;
assign b[57] = 1'b0;
assign a[58] = p3917;
assign b[58] = p3884;
assign a[59] = p3941;
assign b[59] = p3916;
assign a[60] = p3940;
assign b[60] = p3959;
assign a[61] = p3971;
assign b[61] = 1'b0;
assign a[62] = p3977;
assign b[62] = p3970;
assign a[63] = p3972;
assign b[63] = p3974;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[63] = s[63] & p3976;
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
assign o[31] = s[31];
assign o[32] = s[32];
assign o[33] = s[33];
assign o[34] = s[34];
assign o[35] = s[35];
assign o[36] = s[36];
assign o[37] = s[37];
assign o[38] = s[38];
assign o[39] = s[39];
assign o[40] = s[40];
assign o[41] = s[41];
assign o[42] = s[42];
assign o[43] = s[43];
assign o[44] = s[44];
assign o[45] = s[45];
assign o[46] = s[46];
assign o[47] = s[47];
assign o[48] = s[48];
assign o[49] = s[49];
assign o[50] = s[50];
assign o[51] = s[51];
assign o[52] = s[52];
assign o[53] = s[53];
assign o[54] = s[54];
assign o[55] = s[55];
assign o[56] = s[56];
assign o[57] = s[57];
assign o[58] = s[58];
assign o[59] = s[59];
assign o[60] = s[60];
assign o[61] = s[61];
assign o[62] = s[62];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [63:0] a,b;
output [63:0] s;
assign s = a+b;
endmodule
