// 1 2 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 2 1 1 1 1 1 1 1 1 1 2 2 1 1 1 2 2 2 1 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 42 

module main(x,y,o);
input [31:0] x,y;
output [63:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_0_16,ip_0_17,ip_0_18,ip_0_19,ip_0_20,ip_0_21,ip_0_22,ip_0_23,ip_0_24,ip_0_25,ip_0_26,ip_0_27,ip_0_28,ip_0_29,ip_0_30,ip_0_31,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_1_16,ip_1_17,ip_1_18,ip_1_19,ip_1_20,ip_1_21,ip_1_22,ip_1_23,ip_1_24,ip_1_25,ip_1_26,ip_1_27,ip_1_28,ip_1_29,ip_1_30,ip_1_31,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_2_16,ip_2_17,ip_2_18,ip_2_19,ip_2_20,ip_2_21,ip_2_22,ip_2_23,ip_2_24,ip_2_25,ip_2_26,ip_2_27,ip_2_28,ip_2_29,ip_2_30,ip_2_31,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_3_16,ip_3_17,ip_3_18,ip_3_19,ip_3_20,ip_3_21,ip_3_22,ip_3_23,ip_3_24,ip_3_25,ip_3_26,ip_3_27,ip_3_28,ip_3_29,ip_3_30,ip_3_31,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_4_16,ip_4_17,ip_4_18,ip_4_19,ip_4_20,ip_4_21,ip_4_22,ip_4_23,ip_4_24,ip_4_25,ip_4_26,ip_4_27,ip_4_28,ip_4_29,ip_4_30,ip_4_31,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_5_16,ip_5_17,ip_5_18,ip_5_19,ip_5_20,ip_5_21,ip_5_22,ip_5_23,ip_5_24,ip_5_25,ip_5_26,ip_5_27,ip_5_28,ip_5_29,ip_5_30,ip_5_31,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_6_16,ip_6_17,ip_6_18,ip_6_19,ip_6_20,ip_6_21,ip_6_22,ip_6_23,ip_6_24,ip_6_25,ip_6_26,ip_6_27,ip_6_28,ip_6_29,ip_6_30,ip_6_31,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_7_16,ip_7_17,ip_7_18,ip_7_19,ip_7_20,ip_7_21,ip_7_22,ip_7_23,ip_7_24,ip_7_25,ip_7_26,ip_7_27,ip_7_28,ip_7_29,ip_7_30,ip_7_31,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_8_16,ip_8_17,ip_8_18,ip_8_19,ip_8_20,ip_8_21,ip_8_22,ip_8_23,ip_8_24,ip_8_25,ip_8_26,ip_8_27,ip_8_28,ip_8_29,ip_8_30,ip_8_31,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_9_16,ip_9_17,ip_9_18,ip_9_19,ip_9_20,ip_9_21,ip_9_22,ip_9_23,ip_9_24,ip_9_25,ip_9_26,ip_9_27,ip_9_28,ip_9_29,ip_9_30,ip_9_31,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_10_16,ip_10_17,ip_10_18,ip_10_19,ip_10_20,ip_10_21,ip_10_22,ip_10_23,ip_10_24,ip_10_25,ip_10_26,ip_10_27,ip_10_28,ip_10_29,ip_10_30,ip_10_31,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_11_16,ip_11_17,ip_11_18,ip_11_19,ip_11_20,ip_11_21,ip_11_22,ip_11_23,ip_11_24,ip_11_25,ip_11_26,ip_11_27,ip_11_28,ip_11_29,ip_11_30,ip_11_31,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_12_16,ip_12_17,ip_12_18,ip_12_19,ip_12_20,ip_12_21,ip_12_22,ip_12_23,ip_12_24,ip_12_25,ip_12_26,ip_12_27,ip_12_28,ip_12_29,ip_12_30,ip_12_31,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_13_16,ip_13_17,ip_13_18,ip_13_19,ip_13_20,ip_13_21,ip_13_22,ip_13_23,ip_13_24,ip_13_25,ip_13_26,ip_13_27,ip_13_28,ip_13_29,ip_13_30,ip_13_31,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_14_16,ip_14_17,ip_14_18,ip_14_19,ip_14_20,ip_14_21,ip_14_22,ip_14_23,ip_14_24,ip_14_25,ip_14_26,ip_14_27,ip_14_28,ip_14_29,ip_14_30,ip_14_31,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15,ip_15_16,ip_15_17,ip_15_18,ip_15_19,ip_15_20,ip_15_21,ip_15_22,ip_15_23,ip_15_24,ip_15_25,ip_15_26,ip_15_27,ip_15_28,ip_15_29,ip_15_30,ip_15_31,ip_16_0,ip_16_1,ip_16_2,ip_16_3,ip_16_4,ip_16_5,ip_16_6,ip_16_7,ip_16_8,ip_16_9,ip_16_10,ip_16_11,ip_16_12,ip_16_13,ip_16_14,ip_16_15,ip_16_16,ip_16_17,ip_16_18,ip_16_19,ip_16_20,ip_16_21,ip_16_22,ip_16_23,ip_16_24,ip_16_25,ip_16_26,ip_16_27,ip_16_28,ip_16_29,ip_16_30,ip_16_31,ip_17_0,ip_17_1,ip_17_2,ip_17_3,ip_17_4,ip_17_5,ip_17_6,ip_17_7,ip_17_8,ip_17_9,ip_17_10,ip_17_11,ip_17_12,ip_17_13,ip_17_14,ip_17_15,ip_17_16,ip_17_17,ip_17_18,ip_17_19,ip_17_20,ip_17_21,ip_17_22,ip_17_23,ip_17_24,ip_17_25,ip_17_26,ip_17_27,ip_17_28,ip_17_29,ip_17_30,ip_17_31,ip_18_0,ip_18_1,ip_18_2,ip_18_3,ip_18_4,ip_18_5,ip_18_6,ip_18_7,ip_18_8,ip_18_9,ip_18_10,ip_18_11,ip_18_12,ip_18_13,ip_18_14,ip_18_15,ip_18_16,ip_18_17,ip_18_18,ip_18_19,ip_18_20,ip_18_21,ip_18_22,ip_18_23,ip_18_24,ip_18_25,ip_18_26,ip_18_27,ip_18_28,ip_18_29,ip_18_30,ip_18_31,ip_19_0,ip_19_1,ip_19_2,ip_19_3,ip_19_4,ip_19_5,ip_19_6,ip_19_7,ip_19_8,ip_19_9,ip_19_10,ip_19_11,ip_19_12,ip_19_13,ip_19_14,ip_19_15,ip_19_16,ip_19_17,ip_19_18,ip_19_19,ip_19_20,ip_19_21,ip_19_22,ip_19_23,ip_19_24,ip_19_25,ip_19_26,ip_19_27,ip_19_28,ip_19_29,ip_19_30,ip_19_31,ip_20_0,ip_20_1,ip_20_2,ip_20_3,ip_20_4,ip_20_5,ip_20_6,ip_20_7,ip_20_8,ip_20_9,ip_20_10,ip_20_11,ip_20_12,ip_20_13,ip_20_14,ip_20_15,ip_20_16,ip_20_17,ip_20_18,ip_20_19,ip_20_20,ip_20_21,ip_20_22,ip_20_23,ip_20_24,ip_20_25,ip_20_26,ip_20_27,ip_20_28,ip_20_29,ip_20_30,ip_20_31,ip_21_0,ip_21_1,ip_21_2,ip_21_3,ip_21_4,ip_21_5,ip_21_6,ip_21_7,ip_21_8,ip_21_9,ip_21_10,ip_21_11,ip_21_12,ip_21_13,ip_21_14,ip_21_15,ip_21_16,ip_21_17,ip_21_18,ip_21_19,ip_21_20,ip_21_21,ip_21_22,ip_21_23,ip_21_24,ip_21_25,ip_21_26,ip_21_27,ip_21_28,ip_21_29,ip_21_30,ip_21_31,ip_22_0,ip_22_1,ip_22_2,ip_22_3,ip_22_4,ip_22_5,ip_22_6,ip_22_7,ip_22_8,ip_22_9,ip_22_10,ip_22_11,ip_22_12,ip_22_13,ip_22_14,ip_22_15,ip_22_16,ip_22_17,ip_22_18,ip_22_19,ip_22_20,ip_22_21,ip_22_22,ip_22_23,ip_22_24,ip_22_25,ip_22_26,ip_22_27,ip_22_28,ip_22_29,ip_22_30,ip_22_31,ip_23_0,ip_23_1,ip_23_2,ip_23_3,ip_23_4,ip_23_5,ip_23_6,ip_23_7,ip_23_8,ip_23_9,ip_23_10,ip_23_11,ip_23_12,ip_23_13,ip_23_14,ip_23_15,ip_23_16,ip_23_17,ip_23_18,ip_23_19,ip_23_20,ip_23_21,ip_23_22,ip_23_23,ip_23_24,ip_23_25,ip_23_26,ip_23_27,ip_23_28,ip_23_29,ip_23_30,ip_23_31,ip_24_0,ip_24_1,ip_24_2,ip_24_3,ip_24_4,ip_24_5,ip_24_6,ip_24_7,ip_24_8,ip_24_9,ip_24_10,ip_24_11,ip_24_12,ip_24_13,ip_24_14,ip_24_15,ip_24_16,ip_24_17,ip_24_18,ip_24_19,ip_24_20,ip_24_21,ip_24_22,ip_24_23,ip_24_24,ip_24_25,ip_24_26,ip_24_27,ip_24_28,ip_24_29,ip_24_30,ip_24_31,ip_25_0,ip_25_1,ip_25_2,ip_25_3,ip_25_4,ip_25_5,ip_25_6,ip_25_7,ip_25_8,ip_25_9,ip_25_10,ip_25_11,ip_25_12,ip_25_13,ip_25_14,ip_25_15,ip_25_16,ip_25_17,ip_25_18,ip_25_19,ip_25_20,ip_25_21,ip_25_22,ip_25_23,ip_25_24,ip_25_25,ip_25_26,ip_25_27,ip_25_28,ip_25_29,ip_25_30,ip_25_31,ip_26_0,ip_26_1,ip_26_2,ip_26_3,ip_26_4,ip_26_5,ip_26_6,ip_26_7,ip_26_8,ip_26_9,ip_26_10,ip_26_11,ip_26_12,ip_26_13,ip_26_14,ip_26_15,ip_26_16,ip_26_17,ip_26_18,ip_26_19,ip_26_20,ip_26_21,ip_26_22,ip_26_23,ip_26_24,ip_26_25,ip_26_26,ip_26_27,ip_26_28,ip_26_29,ip_26_30,ip_26_31,ip_27_0,ip_27_1,ip_27_2,ip_27_3,ip_27_4,ip_27_5,ip_27_6,ip_27_7,ip_27_8,ip_27_9,ip_27_10,ip_27_11,ip_27_12,ip_27_13,ip_27_14,ip_27_15,ip_27_16,ip_27_17,ip_27_18,ip_27_19,ip_27_20,ip_27_21,ip_27_22,ip_27_23,ip_27_24,ip_27_25,ip_27_26,ip_27_27,ip_27_28,ip_27_29,ip_27_30,ip_27_31,ip_28_0,ip_28_1,ip_28_2,ip_28_3,ip_28_4,ip_28_5,ip_28_6,ip_28_7,ip_28_8,ip_28_9,ip_28_10,ip_28_11,ip_28_12,ip_28_13,ip_28_14,ip_28_15,ip_28_16,ip_28_17,ip_28_18,ip_28_19,ip_28_20,ip_28_21,ip_28_22,ip_28_23,ip_28_24,ip_28_25,ip_28_26,ip_28_27,ip_28_28,ip_28_29,ip_28_30,ip_28_31,ip_29_0,ip_29_1,ip_29_2,ip_29_3,ip_29_4,ip_29_5,ip_29_6,ip_29_7,ip_29_8,ip_29_9,ip_29_10,ip_29_11,ip_29_12,ip_29_13,ip_29_14,ip_29_15,ip_29_16,ip_29_17,ip_29_18,ip_29_19,ip_29_20,ip_29_21,ip_29_22,ip_29_23,ip_29_24,ip_29_25,ip_29_26,ip_29_27,ip_29_28,ip_29_29,ip_29_30,ip_29_31,ip_30_0,ip_30_1,ip_30_2,ip_30_3,ip_30_4,ip_30_5,ip_30_6,ip_30_7,ip_30_8,ip_30_9,ip_30_10,ip_30_11,ip_30_12,ip_30_13,ip_30_14,ip_30_15,ip_30_16,ip_30_17,ip_30_18,ip_30_19,ip_30_20,ip_30_21,ip_30_22,ip_30_23,ip_30_24,ip_30_25,ip_30_26,ip_30_27,ip_30_28,ip_30_29,ip_30_30,ip_30_31,ip_31_0,ip_31_1,ip_31_2,ip_31_3,ip_31_4,ip_31_5,ip_31_6,ip_31_7,ip_31_8,ip_31_9,ip_31_10,ip_31_11,ip_31_12,ip_31_13,ip_31_14,ip_31_15,ip_31_16,ip_31_17,ip_31_18,ip_31_19,ip_31_20,ip_31_21,ip_31_22,ip_31_23,ip_31_24,ip_31_25,ip_31_26,ip_31_27,ip_31_28,ip_31_29,ip_31_30,ip_31_31;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149,p1150,p1151,p1152,p1153,p1154,p1155,p1156,p1157,p1158,p1159,p1160,p1161,p1162,p1163,p1164,p1165,p1166,p1167,p1168,p1169,p1170,p1171,p1172,p1173,p1174,p1175,p1176,p1177,p1178,p1179,p1180,p1181,p1182,p1183,p1184,p1185,p1186,p1187,p1188,p1189,p1190,p1191,p1192,p1193,p1194,p1195,p1196,p1197,p1198,p1199,p1200,p1201,p1202,p1203,p1204,p1205,p1206,p1207,p1208,p1209,p1210,p1211,p1212,p1213,p1214,p1215,p1216,p1217,p1218,p1219,p1220,p1221,p1222,p1223,p1224,p1225,p1226,p1227,p1228,p1229,p1230,p1231,p1232,p1233,p1234,p1235,p1236,p1237,p1238,p1239,p1240,p1241,p1242,p1243,p1244,p1245,p1246,p1247,p1248,p1249,p1250,p1251,p1252,p1253,p1254,p1255,p1256,p1257,p1258,p1259,p1260,p1261,p1262,p1263,p1264,p1265,p1266,p1267,p1268,p1269,p1270,p1271,p1272,p1273,p1274,p1275,p1276,p1277,p1278,p1279,p1280,p1281,p1282,p1283,p1284,p1285,p1286,p1287,p1288,p1289,p1290,p1291,p1292,p1293,p1294,p1295,p1296,p1297,p1298,p1299,p1300,p1301,p1302,p1303,p1304,p1305,p1306,p1307,p1308,p1309,p1310,p1311,p1312,p1313,p1314,p1315,p1316,p1317,p1318,p1319,p1320,p1321,p1322,p1323,p1324,p1325,p1326,p1327,p1328,p1329,p1330,p1331,p1332,p1333,p1334,p1335,p1336,p1337,p1338,p1339,p1340,p1341,p1342,p1343,p1344,p1345,p1346,p1347,p1348,p1349,p1350,p1351,p1352,p1353,p1354,p1355,p1356,p1357,p1358,p1359,p1360,p1361,p1362,p1363,p1364,p1365,p1366,p1367,p1368,p1369,p1370,p1371,p1372,p1373,p1374,p1375,p1376,p1377,p1378,p1379,p1380,p1381,p1382,p1383,p1384,p1385,p1386,p1387,p1388,p1389,p1390,p1391,p1392,p1393,p1394,p1395,p1396,p1397,p1398,p1399,p1400,p1401,p1402,p1403,p1404,p1405,p1406,p1407,p1408,p1409,p1410,p1411,p1412,p1413,p1414,p1415,p1416,p1417,p1418,p1419,p1420,p1421,p1422,p1423,p1424,p1425,p1426,p1427,p1428,p1429,p1430,p1431,p1432,p1433,p1434,p1435,p1436,p1437,p1438,p1439,p1440,p1441,p1442,p1443,p1444,p1445,p1446,p1447,p1448,p1449,p1450,p1451,p1452,p1453,p1454,p1455,p1456,p1457,p1458,p1459,p1460,p1461,p1462,p1463,p1464,p1465,p1466,p1467,p1468,p1469,p1470,p1471,p1472,p1473,p1474,p1475,p1476,p1477,p1478,p1479,p1480,p1481,p1482,p1483,p1484,p1485,p1486,p1487,p1488,p1489,p1490,p1491,p1492,p1493,p1494,p1495,p1496,p1497,p1498,p1499,p1500,p1501,p1502,p1503,p1504,p1505,p1506,p1507,p1508,p1509,p1510,p1511,p1512,p1513,p1514,p1515,p1516,p1517,p1518,p1519,p1520,p1521,p1522,p1523,p1524,p1525,p1526,p1527,p1528,p1529,p1530,p1531,p1532,p1533,p1534,p1535,p1536,p1537,p1538,p1539,p1540,p1541,p1542,p1543,p1544,p1545,p1546,p1547,p1548,p1549,p1550,p1551,p1552,p1553,p1554,p1555,p1556,p1557,p1558,p1559,p1560,p1561,p1562,p1563,p1564,p1565,p1566,p1567,p1568,p1569,p1570,p1571,p1572,p1573,p1574,p1575,p1576,p1577,p1578,p1579,p1580,p1581,p1582,p1583,p1584,p1585,p1586,p1587,p1588,p1589,p1590,p1591,p1592,p1593,p1594,p1595,p1596,p1597,p1598,p1599,p1600,p1601,p1602,p1603,p1604,p1605,p1606,p1607,p1608,p1609,p1610,p1611,p1612,p1613,p1614,p1615,p1616,p1617,p1618,p1619,p1620,p1621,p1622,p1623,p1624,p1625,p1626,p1627,p1628,p1629,p1630,p1631,p1632,p1633,p1634,p1635,p1636,p1637,p1638,p1639,p1640,p1641,p1642,p1643,p1644,p1645,p1646,p1647,p1648,p1649,p1650,p1651,p1652,p1653,p1654,p1655,p1656,p1657,p1658,p1659,p1660,p1661,p1662,p1663,p1664,p1665,p1666,p1667,p1668,p1669,p1670,p1671,p1672,p1673,p1674,p1675,p1676,p1677,p1678,p1679,p1680,p1681,p1682,p1683,p1684,p1685,p1686,p1687,p1688,p1689,p1690,p1691,p1692,p1693,p1694,p1695,p1696,p1697,p1698,p1699,p1700,p1701,p1702,p1703,p1704,p1705,p1706,p1707,p1708,p1709,p1710,p1711,p1712,p1713,p1714,p1715,p1716,p1717,p1718,p1719,p1720,p1721,p1722,p1723,p1724,p1725,p1726,p1727,p1728,p1729,p1730,p1731,p1732,p1733,p1734,p1735,p1736,p1737,p1738,p1739,p1740,p1741,p1742,p1743,p1744,p1745,p1746,p1747,p1748,p1749,p1750,p1751,p1752,p1753,p1754,p1755,p1756,p1757,p1758,p1759,p1760,p1761,p1762,p1763,p1764,p1765,p1766,p1767,p1768,p1769,p1770,p1771,p1772,p1773,p1774,p1775,p1776,p1777,p1778,p1779,p1780,p1781,p1782,p1783,p1784,p1785,p1786,p1787,p1788,p1789,p1790,p1791,p1792,p1793,p1794,p1795,p1796,p1797,p1798,p1799,p1800,p1801,p1802,p1803,p1804,p1805,p1806,p1807,p1808,p1809,p1810,p1811,p1812,p1813,p1814,p1815,p1816,p1817,p1818,p1819,p1820,p1821,p1822,p1823,p1824,p1825,p1826,p1827,p1828,p1829,p1830,p1831,p1832,p1833,p1834,p1835,p1836,p1837,p1838,p1839,p1840,p1841,p1842,p1843,p1844,p1845,p1846,p1847,p1848,p1849,p1850,p1851,p1852,p1853,p1854,p1855,p1856,p1857,p1858,p1859,p1860,p1861,p1862,p1863,p1864,p1865,p1866,p1867,p1868,p1869,p1870,p1871,p1872,p1873,p1874,p1875,p1876,p1877,p1878,p1879,p1880,p1881,p1882,p1883,p1884,p1885,p1886,p1887,p1888,p1889,p1890,p1891,p1892,p1893,p1894,p1895,p1896,p1897,p1898,p1899,p1900,p1901,p1902,p1903,p1904,p1905,p1906,p1907,p1908,p1909,p1910,p1911,p1912,p1913,p1914,p1915,p1916,p1917,p1918,p1919,p1920,p1921,p1922,p1923,p1924,p1925,p1926,p1927,p1928,p1929,p1930,p1931,p1932,p1933,p1934,p1935,p1936,p1937,p1938,p1939,p1940,p1941,p1942,p1943,p1944,p1945,p1946,p1947,p1948,p1949,p1950,p1951,p1952,p1953,p1954,p1955,p1956,p1957,p1958,p1959,p1960,p1961,p1962,p1963,p1964,p1965,p1966,p1967,p1968,p1969,p1970,p1971,p1972,p1973,p1974,p1975,p1976,p1977,p1978,p1979,p1980,p1981,p1982,p1983,p1984,p1985,p1986,p1987,p1988,p1989,p1990,p1991,p1992,p1993,p1994,p1995,p1996,p1997,p1998,p1999,p2000,p2001,p2002,p2003,p2004,p2005,p2006,p2007,p2008,p2009,p2010,p2011,p2012,p2013,p2014,p2015,p2016,p2017,p2018,p2019,p2020,p2021,p2022,p2023,p2024,p2025,p2026,p2027,p2028,p2029,p2030,p2031,p2032,p2033,p2034,p2035,p2036,p2037,p2038,p2039,p2040,p2041,p2042,p2043,p2044,p2045,p2046,p2047,p2048,p2049,p2050,p2051,p2052,p2053,p2054,p2055,p2056,p2057,p2058,p2059,p2060,p2061,p2062,p2063,p2064,p2065,p2066,p2067,p2068,p2069,p2070,p2071,p2072,p2073,p2074,p2075,p2076,p2077,p2078,p2079,p2080,p2081,p2082,p2083,p2084,p2085,p2086,p2087,p2088,p2089,p2090,p2091,p2092,p2093,p2094,p2095,p2096,p2097,p2098,p2099,p2100,p2101,p2102,p2103,p2104,p2105,p2106,p2107,p2108,p2109,p2110,p2111,p2112,p2113,p2114,p2115,p2116,p2117,p2118,p2119,p2120,p2121,p2122,p2123,p2124,p2125,p2126,p2127,p2128,p2129,p2130,p2131,p2132,p2133,p2134,p2135,p2136,p2137,p2138,p2139,p2140,p2141,p2142,p2143,p2144,p2145,p2146,p2147,p2148,p2149,p2150,p2151,p2152,p2153,p2154,p2155,p2156,p2157,p2158,p2159,p2160,p2161,p2162,p2163,p2164,p2165,p2166,p2167,p2168,p2169,p2170,p2171,p2172,p2173,p2174,p2175,p2176,p2177,p2178,p2179,p2180,p2181,p2182,p2183,p2184,p2185,p2186,p2187,p2188,p2189,p2190,p2191,p2192,p2193,p2194,p2195,p2196,p2197,p2198,p2199,p2200,p2201,p2202,p2203,p2204,p2205,p2206,p2207,p2208,p2209,p2210,p2211,p2212,p2213,p2214,p2215,p2216,p2217,p2218,p2219,p2220,p2221,p2222,p2223,p2224,p2225,p2226,p2227,p2228,p2229,p2230,p2231,p2232,p2233,p2234,p2235,p2236,p2237,p2238,p2239,p2240,p2241,p2242,p2243,p2244,p2245,p2246,p2247,p2248,p2249,p2250,p2251,p2252,p2253,p2254,p2255,p2256,p2257,p2258,p2259,p2260,p2261,p2262,p2263,p2264,p2265,p2266,p2267,p2268,p2269,p2270,p2271,p2272,p2273,p2274,p2275,p2276,p2277,p2278,p2279,p2280,p2281,p2282,p2283,p2284,p2285,p2286,p2287,p2288,p2289,p2290,p2291,p2292,p2293,p2294,p2295,p2296,p2297,p2298,p2299,p2300,p2301,p2302,p2303,p2304,p2305,p2306,p2307,p2308,p2309,p2310,p2311,p2312,p2313,p2314,p2315,p2316,p2317,p2318,p2319,p2320,p2321,p2322,p2323,p2324,p2325,p2326,p2327,p2328,p2329,p2330,p2331,p2332,p2333,p2334,p2335,p2336,p2337,p2338,p2339,p2340,p2341,p2342,p2343,p2344,p2345,p2346,p2347,p2348,p2349,p2350,p2351,p2352,p2353,p2354,p2355,p2356,p2357,p2358,p2359,p2360,p2361,p2362,p2363,p2364,p2365,p2366,p2367,p2368,p2369,p2370,p2371,p2372,p2373,p2374,p2375,p2376,p2377,p2378,p2379,p2380,p2381,p2382,p2383,p2384,p2385,p2386,p2387,p2388,p2389,p2390,p2391,p2392,p2393,p2394,p2395,p2396,p2397,p2398,p2399,p2400,p2401,p2402,p2403,p2404,p2405,p2406,p2407,p2408,p2409,p2410,p2411,p2412,p2413,p2414,p2415,p2416,p2417,p2418,p2419,p2420,p2421,p2422,p2423,p2424,p2425,p2426,p2427,p2428,p2429,p2430,p2431,p2432,p2433,p2434,p2435,p2436,p2437,p2438,p2439,p2440,p2441,p2442,p2443,p2444,p2445,p2446,p2447,p2448,p2449,p2450,p2451,p2452,p2453,p2454,p2455,p2456,p2457,p2458,p2459,p2460,p2461,p2462,p2463,p2464,p2465,p2466,p2467,p2468,p2469,p2470,p2471,p2472,p2473,p2474,p2475,p2476,p2477,p2478,p2479,p2480,p2481,p2482,p2483,p2484,p2485,p2486,p2487,p2488,p2489,p2490,p2491,p2492,p2493,p2494,p2495,p2496,p2497,p2498,p2499,p2500,p2501,p2502,p2503,p2504,p2505,p2506,p2507,p2508,p2509,p2510,p2511,p2512,p2513,p2514,p2515,p2516,p2517,p2518,p2519,p2520,p2521,p2522,p2523,p2524,p2525,p2526,p2527,p2528,p2529,p2530,p2531,p2532,p2533,p2534,p2535,p2536,p2537,p2538,p2539,p2540,p2541,p2542,p2543,p2544,p2545,p2546,p2547,p2548,p2549,p2550,p2551,p2552,p2553,p2554,p2555,p2556,p2557,p2558,p2559,p2560,p2561,p2562,p2563,p2564,p2565,p2566,p2567,p2568,p2569,p2570,p2571,p2572,p2573,p2574,p2575,p2576,p2577,p2578,p2579,p2580,p2581,p2582,p2583,p2584,p2585,p2586,p2587,p2588,p2589,p2590,p2591,p2592,p2593,p2594,p2595,p2596,p2597,p2598,p2599,p2600,p2601,p2602,p2603,p2604,p2605,p2606,p2607,p2608,p2609,p2610,p2611,p2612,p2613,p2614,p2615,p2616,p2617,p2618,p2619,p2620,p2621,p2622,p2623,p2624,p2625,p2626,p2627,p2628,p2629,p2630,p2631,p2632,p2633,p2634,p2635,p2636,p2637,p2638,p2639,p2640,p2641,p2642,p2643,p2644,p2645,p2646,p2647,p2648,p2649,p2650,p2651,p2652,p2653,p2654,p2655,p2656,p2657,p2658,p2659,p2660,p2661,p2662,p2663,p2664,p2665,p2666,p2667,p2668,p2669,p2670,p2671,p2672,p2673,p2674,p2675,p2676,p2677,p2678,p2679,p2680,p2681,p2682,p2683,p2684,p2685,p2686,p2687,p2688,p2689,p2690,p2691,p2692,p2693,p2694,p2695,p2696,p2697,p2698,p2699,p2700,p2701,p2702,p2703,p2704,p2705,p2706,p2707,p2708,p2709,p2710,p2711,p2712,p2713,p2714,p2715,p2716,p2717,p2718,p2719,p2720,p2721,p2722,p2723,p2724,p2725,p2726,p2727,p2728,p2729,p2730,p2731,p2732,p2733,p2734,p2735,p2736,p2737,p2738,p2739,p2740,p2741,p2742,p2743,p2744,p2745,p2746,p2747,p2748,p2749,p2750,p2751,p2752,p2753,p2754,p2755,p2756,p2757,p2758,p2759,p2760,p2761,p2762,p2763,p2764,p2765,p2766,p2767,p2768,p2769,p2770,p2771,p2772,p2773,p2774,p2775,p2776,p2777,p2778,p2779,p2780,p2781,p2782,p2783,p2784,p2785,p2786,p2787,p2788,p2789,p2790,p2791,p2792,p2793,p2794,p2795,p2796,p2797,p2798,p2799,p2800,p2801,p2802,p2803,p2804,p2805,p2806,p2807,p2808,p2809,p2810,p2811,p2812,p2813,p2814,p2815,p2816,p2817,p2818,p2819,p2820,p2821,p2822,p2823,p2824,p2825,p2826,p2827,p2828,p2829,p2830,p2831,p2832,p2833,p2834,p2835,p2836,p2837,p2838,p2839,p2840,p2841,p2842,p2843,p2844,p2845,p2846,p2847,p2848,p2849,p2850,p2851,p2852,p2853,p2854,p2855,p2856,p2857,p2858,p2859,p2860,p2861,p2862,p2863,p2864,p2865,p2866,p2867,p2868,p2869,p2870,p2871,p2872,p2873,p2874,p2875,p2876,p2877,p2878,p2879;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_0_16,x[0],y[16]);
and and17(ip_0_17,x[0],y[17]);
and and18(ip_0_18,x[0],y[18]);
and and19(ip_0_19,x[0],y[19]);
and and20(ip_0_20,x[0],y[20]);
and and21(ip_0_21,x[0],y[21]);
and and22(ip_0_22,x[0],y[22]);
and and23(ip_0_23,x[0],y[23]);
and and24(ip_0_24,x[0],y[24]);
and and25(ip_0_25,x[0],y[25]);
and and26(ip_0_26,x[0],y[26]);
and and27(ip_0_27,x[0],y[27]);
and and28(ip_0_28,x[0],y[28]);
and and29(ip_0_29,x[0],y[29]);
and and30(ip_0_30,x[0],y[30]);
and and31(ip_0_31,x[0],y[31]);
and and32(ip_1_0,x[1],y[0]);
and and33(ip_1_1,x[1],y[1]);
and and34(ip_1_2,x[1],y[2]);
and and35(ip_1_3,x[1],y[3]);
and and36(ip_1_4,x[1],y[4]);
and and37(ip_1_5,x[1],y[5]);
and and38(ip_1_6,x[1],y[6]);
and and39(ip_1_7,x[1],y[7]);
and and40(ip_1_8,x[1],y[8]);
and and41(ip_1_9,x[1],y[9]);
and and42(ip_1_10,x[1],y[10]);
and and43(ip_1_11,x[1],y[11]);
and and44(ip_1_12,x[1],y[12]);
and and45(ip_1_13,x[1],y[13]);
and and46(ip_1_14,x[1],y[14]);
and and47(ip_1_15,x[1],y[15]);
and and48(ip_1_16,x[1],y[16]);
and and49(ip_1_17,x[1],y[17]);
and and50(ip_1_18,x[1],y[18]);
and and51(ip_1_19,x[1],y[19]);
and and52(ip_1_20,x[1],y[20]);
and and53(ip_1_21,x[1],y[21]);
and and54(ip_1_22,x[1],y[22]);
and and55(ip_1_23,x[1],y[23]);
and and56(ip_1_24,x[1],y[24]);
and and57(ip_1_25,x[1],y[25]);
and and58(ip_1_26,x[1],y[26]);
and and59(ip_1_27,x[1],y[27]);
and and60(ip_1_28,x[1],y[28]);
and and61(ip_1_29,x[1],y[29]);
and and62(ip_1_30,x[1],y[30]);
and and63(ip_1_31,x[1],y[31]);
and and64(ip_2_0,x[2],y[0]);
and and65(ip_2_1,x[2],y[1]);
and and66(ip_2_2,x[2],y[2]);
and and67(ip_2_3,x[2],y[3]);
and and68(ip_2_4,x[2],y[4]);
and and69(ip_2_5,x[2],y[5]);
and and70(ip_2_6,x[2],y[6]);
and and71(ip_2_7,x[2],y[7]);
and and72(ip_2_8,x[2],y[8]);
and and73(ip_2_9,x[2],y[9]);
and and74(ip_2_10,x[2],y[10]);
and and75(ip_2_11,x[2],y[11]);
and and76(ip_2_12,x[2],y[12]);
and and77(ip_2_13,x[2],y[13]);
and and78(ip_2_14,x[2],y[14]);
and and79(ip_2_15,x[2],y[15]);
and and80(ip_2_16,x[2],y[16]);
and and81(ip_2_17,x[2],y[17]);
and and82(ip_2_18,x[2],y[18]);
and and83(ip_2_19,x[2],y[19]);
and and84(ip_2_20,x[2],y[20]);
and and85(ip_2_21,x[2],y[21]);
and and86(ip_2_22,x[2],y[22]);
and and87(ip_2_23,x[2],y[23]);
and and88(ip_2_24,x[2],y[24]);
and and89(ip_2_25,x[2],y[25]);
and and90(ip_2_26,x[2],y[26]);
and and91(ip_2_27,x[2],y[27]);
and and92(ip_2_28,x[2],y[28]);
and and93(ip_2_29,x[2],y[29]);
and and94(ip_2_30,x[2],y[30]);
and and95(ip_2_31,x[2],y[31]);
and and96(ip_3_0,x[3],y[0]);
and and97(ip_3_1,x[3],y[1]);
and and98(ip_3_2,x[3],y[2]);
and and99(ip_3_3,x[3],y[3]);
and and100(ip_3_4,x[3],y[4]);
and and101(ip_3_5,x[3],y[5]);
and and102(ip_3_6,x[3],y[6]);
and and103(ip_3_7,x[3],y[7]);
and and104(ip_3_8,x[3],y[8]);
and and105(ip_3_9,x[3],y[9]);
and and106(ip_3_10,x[3],y[10]);
and and107(ip_3_11,x[3],y[11]);
and and108(ip_3_12,x[3],y[12]);
and and109(ip_3_13,x[3],y[13]);
and and110(ip_3_14,x[3],y[14]);
and and111(ip_3_15,x[3],y[15]);
and and112(ip_3_16,x[3],y[16]);
and and113(ip_3_17,x[3],y[17]);
and and114(ip_3_18,x[3],y[18]);
and and115(ip_3_19,x[3],y[19]);
and and116(ip_3_20,x[3],y[20]);
and and117(ip_3_21,x[3],y[21]);
and and118(ip_3_22,x[3],y[22]);
and and119(ip_3_23,x[3],y[23]);
and and120(ip_3_24,x[3],y[24]);
and and121(ip_3_25,x[3],y[25]);
and and122(ip_3_26,x[3],y[26]);
and and123(ip_3_27,x[3],y[27]);
and and124(ip_3_28,x[3],y[28]);
and and125(ip_3_29,x[3],y[29]);
and and126(ip_3_30,x[3],y[30]);
and and127(ip_3_31,x[3],y[31]);
and and128(ip_4_0,x[4],y[0]);
and and129(ip_4_1,x[4],y[1]);
and and130(ip_4_2,x[4],y[2]);
and and131(ip_4_3,x[4],y[3]);
and and132(ip_4_4,x[4],y[4]);
and and133(ip_4_5,x[4],y[5]);
and and134(ip_4_6,x[4],y[6]);
and and135(ip_4_7,x[4],y[7]);
and and136(ip_4_8,x[4],y[8]);
and and137(ip_4_9,x[4],y[9]);
and and138(ip_4_10,x[4],y[10]);
and and139(ip_4_11,x[4],y[11]);
and and140(ip_4_12,x[4],y[12]);
and and141(ip_4_13,x[4],y[13]);
and and142(ip_4_14,x[4],y[14]);
and and143(ip_4_15,x[4],y[15]);
and and144(ip_4_16,x[4],y[16]);
and and145(ip_4_17,x[4],y[17]);
and and146(ip_4_18,x[4],y[18]);
and and147(ip_4_19,x[4],y[19]);
and and148(ip_4_20,x[4],y[20]);
and and149(ip_4_21,x[4],y[21]);
and and150(ip_4_22,x[4],y[22]);
and and151(ip_4_23,x[4],y[23]);
and and152(ip_4_24,x[4],y[24]);
and and153(ip_4_25,x[4],y[25]);
and and154(ip_4_26,x[4],y[26]);
and and155(ip_4_27,x[4],y[27]);
and and156(ip_4_28,x[4],y[28]);
and and157(ip_4_29,x[4],y[29]);
and and158(ip_4_30,x[4],y[30]);
and and159(ip_4_31,x[4],y[31]);
and and160(ip_5_0,x[5],y[0]);
and and161(ip_5_1,x[5],y[1]);
and and162(ip_5_2,x[5],y[2]);
and and163(ip_5_3,x[5],y[3]);
and and164(ip_5_4,x[5],y[4]);
and and165(ip_5_5,x[5],y[5]);
and and166(ip_5_6,x[5],y[6]);
and and167(ip_5_7,x[5],y[7]);
and and168(ip_5_8,x[5],y[8]);
and and169(ip_5_9,x[5],y[9]);
and and170(ip_5_10,x[5],y[10]);
and and171(ip_5_11,x[5],y[11]);
and and172(ip_5_12,x[5],y[12]);
and and173(ip_5_13,x[5],y[13]);
and and174(ip_5_14,x[5],y[14]);
and and175(ip_5_15,x[5],y[15]);
and and176(ip_5_16,x[5],y[16]);
and and177(ip_5_17,x[5],y[17]);
and and178(ip_5_18,x[5],y[18]);
and and179(ip_5_19,x[5],y[19]);
and and180(ip_5_20,x[5],y[20]);
and and181(ip_5_21,x[5],y[21]);
and and182(ip_5_22,x[5],y[22]);
and and183(ip_5_23,x[5],y[23]);
and and184(ip_5_24,x[5],y[24]);
and and185(ip_5_25,x[5],y[25]);
and and186(ip_5_26,x[5],y[26]);
and and187(ip_5_27,x[5],y[27]);
and and188(ip_5_28,x[5],y[28]);
and and189(ip_5_29,x[5],y[29]);
and and190(ip_5_30,x[5],y[30]);
and and191(ip_5_31,x[5],y[31]);
and and192(ip_6_0,x[6],y[0]);
and and193(ip_6_1,x[6],y[1]);
and and194(ip_6_2,x[6],y[2]);
and and195(ip_6_3,x[6],y[3]);
and and196(ip_6_4,x[6],y[4]);
and and197(ip_6_5,x[6],y[5]);
and and198(ip_6_6,x[6],y[6]);
and and199(ip_6_7,x[6],y[7]);
and and200(ip_6_8,x[6],y[8]);
and and201(ip_6_9,x[6],y[9]);
and and202(ip_6_10,x[6],y[10]);
and and203(ip_6_11,x[6],y[11]);
and and204(ip_6_12,x[6],y[12]);
and and205(ip_6_13,x[6],y[13]);
and and206(ip_6_14,x[6],y[14]);
and and207(ip_6_15,x[6],y[15]);
and and208(ip_6_16,x[6],y[16]);
and and209(ip_6_17,x[6],y[17]);
and and210(ip_6_18,x[6],y[18]);
and and211(ip_6_19,x[6],y[19]);
and and212(ip_6_20,x[6],y[20]);
and and213(ip_6_21,x[6],y[21]);
and and214(ip_6_22,x[6],y[22]);
and and215(ip_6_23,x[6],y[23]);
and and216(ip_6_24,x[6],y[24]);
and and217(ip_6_25,x[6],y[25]);
and and218(ip_6_26,x[6],y[26]);
and and219(ip_6_27,x[6],y[27]);
and and220(ip_6_28,x[6],y[28]);
and and221(ip_6_29,x[6],y[29]);
and and222(ip_6_30,x[6],y[30]);
and and223(ip_6_31,x[6],y[31]);
and and224(ip_7_0,x[7],y[0]);
and and225(ip_7_1,x[7],y[1]);
and and226(ip_7_2,x[7],y[2]);
and and227(ip_7_3,x[7],y[3]);
and and228(ip_7_4,x[7],y[4]);
and and229(ip_7_5,x[7],y[5]);
and and230(ip_7_6,x[7],y[6]);
and and231(ip_7_7,x[7],y[7]);
and and232(ip_7_8,x[7],y[8]);
and and233(ip_7_9,x[7],y[9]);
and and234(ip_7_10,x[7],y[10]);
and and235(ip_7_11,x[7],y[11]);
and and236(ip_7_12,x[7],y[12]);
and and237(ip_7_13,x[7],y[13]);
and and238(ip_7_14,x[7],y[14]);
and and239(ip_7_15,x[7],y[15]);
and and240(ip_7_16,x[7],y[16]);
and and241(ip_7_17,x[7],y[17]);
and and242(ip_7_18,x[7],y[18]);
and and243(ip_7_19,x[7],y[19]);
and and244(ip_7_20,x[7],y[20]);
and and245(ip_7_21,x[7],y[21]);
and and246(ip_7_22,x[7],y[22]);
and and247(ip_7_23,x[7],y[23]);
and and248(ip_7_24,x[7],y[24]);
and and249(ip_7_25,x[7],y[25]);
and and250(ip_7_26,x[7],y[26]);
and and251(ip_7_27,x[7],y[27]);
and and252(ip_7_28,x[7],y[28]);
and and253(ip_7_29,x[7],y[29]);
and and254(ip_7_30,x[7],y[30]);
and and255(ip_7_31,x[7],y[31]);
and and256(ip_8_0,x[8],y[0]);
and and257(ip_8_1,x[8],y[1]);
and and258(ip_8_2,x[8],y[2]);
and and259(ip_8_3,x[8],y[3]);
and and260(ip_8_4,x[8],y[4]);
and and261(ip_8_5,x[8],y[5]);
and and262(ip_8_6,x[8],y[6]);
and and263(ip_8_7,x[8],y[7]);
and and264(ip_8_8,x[8],y[8]);
and and265(ip_8_9,x[8],y[9]);
and and266(ip_8_10,x[8],y[10]);
and and267(ip_8_11,x[8],y[11]);
and and268(ip_8_12,x[8],y[12]);
and and269(ip_8_13,x[8],y[13]);
and and270(ip_8_14,x[8],y[14]);
and and271(ip_8_15,x[8],y[15]);
and and272(ip_8_16,x[8],y[16]);
and and273(ip_8_17,x[8],y[17]);
and and274(ip_8_18,x[8],y[18]);
and and275(ip_8_19,x[8],y[19]);
and and276(ip_8_20,x[8],y[20]);
and and277(ip_8_21,x[8],y[21]);
and and278(ip_8_22,x[8],y[22]);
and and279(ip_8_23,x[8],y[23]);
and and280(ip_8_24,x[8],y[24]);
and and281(ip_8_25,x[8],y[25]);
and and282(ip_8_26,x[8],y[26]);
and and283(ip_8_27,x[8],y[27]);
and and284(ip_8_28,x[8],y[28]);
and and285(ip_8_29,x[8],y[29]);
and and286(ip_8_30,x[8],y[30]);
and and287(ip_8_31,x[8],y[31]);
and and288(ip_9_0,x[9],y[0]);
and and289(ip_9_1,x[9],y[1]);
and and290(ip_9_2,x[9],y[2]);
and and291(ip_9_3,x[9],y[3]);
and and292(ip_9_4,x[9],y[4]);
and and293(ip_9_5,x[9],y[5]);
and and294(ip_9_6,x[9],y[6]);
and and295(ip_9_7,x[9],y[7]);
and and296(ip_9_8,x[9],y[8]);
and and297(ip_9_9,x[9],y[9]);
and and298(ip_9_10,x[9],y[10]);
and and299(ip_9_11,x[9],y[11]);
and and300(ip_9_12,x[9],y[12]);
and and301(ip_9_13,x[9],y[13]);
and and302(ip_9_14,x[9],y[14]);
and and303(ip_9_15,x[9],y[15]);
and and304(ip_9_16,x[9],y[16]);
and and305(ip_9_17,x[9],y[17]);
and and306(ip_9_18,x[9],y[18]);
and and307(ip_9_19,x[9],y[19]);
and and308(ip_9_20,x[9],y[20]);
and and309(ip_9_21,x[9],y[21]);
and and310(ip_9_22,x[9],y[22]);
and and311(ip_9_23,x[9],y[23]);
and and312(ip_9_24,x[9],y[24]);
and and313(ip_9_25,x[9],y[25]);
and and314(ip_9_26,x[9],y[26]);
and and315(ip_9_27,x[9],y[27]);
and and316(ip_9_28,x[9],y[28]);
and and317(ip_9_29,x[9],y[29]);
and and318(ip_9_30,x[9],y[30]);
and and319(ip_9_31,x[9],y[31]);
and and320(ip_10_0,x[10],y[0]);
and and321(ip_10_1,x[10],y[1]);
and and322(ip_10_2,x[10],y[2]);
and and323(ip_10_3,x[10],y[3]);
and and324(ip_10_4,x[10],y[4]);
and and325(ip_10_5,x[10],y[5]);
and and326(ip_10_6,x[10],y[6]);
and and327(ip_10_7,x[10],y[7]);
and and328(ip_10_8,x[10],y[8]);
and and329(ip_10_9,x[10],y[9]);
and and330(ip_10_10,x[10],y[10]);
and and331(ip_10_11,x[10],y[11]);
and and332(ip_10_12,x[10],y[12]);
and and333(ip_10_13,x[10],y[13]);
and and334(ip_10_14,x[10],y[14]);
and and335(ip_10_15,x[10],y[15]);
and and336(ip_10_16,x[10],y[16]);
and and337(ip_10_17,x[10],y[17]);
and and338(ip_10_18,x[10],y[18]);
and and339(ip_10_19,x[10],y[19]);
and and340(ip_10_20,x[10],y[20]);
and and341(ip_10_21,x[10],y[21]);
and and342(ip_10_22,x[10],y[22]);
and and343(ip_10_23,x[10],y[23]);
and and344(ip_10_24,x[10],y[24]);
and and345(ip_10_25,x[10],y[25]);
and and346(ip_10_26,x[10],y[26]);
and and347(ip_10_27,x[10],y[27]);
and and348(ip_10_28,x[10],y[28]);
and and349(ip_10_29,x[10],y[29]);
and and350(ip_10_30,x[10],y[30]);
and and351(ip_10_31,x[10],y[31]);
and and352(ip_11_0,x[11],y[0]);
and and353(ip_11_1,x[11],y[1]);
and and354(ip_11_2,x[11],y[2]);
and and355(ip_11_3,x[11],y[3]);
and and356(ip_11_4,x[11],y[4]);
and and357(ip_11_5,x[11],y[5]);
and and358(ip_11_6,x[11],y[6]);
and and359(ip_11_7,x[11],y[7]);
and and360(ip_11_8,x[11],y[8]);
and and361(ip_11_9,x[11],y[9]);
and and362(ip_11_10,x[11],y[10]);
and and363(ip_11_11,x[11],y[11]);
and and364(ip_11_12,x[11],y[12]);
and and365(ip_11_13,x[11],y[13]);
and and366(ip_11_14,x[11],y[14]);
and and367(ip_11_15,x[11],y[15]);
and and368(ip_11_16,x[11],y[16]);
and and369(ip_11_17,x[11],y[17]);
and and370(ip_11_18,x[11],y[18]);
and and371(ip_11_19,x[11],y[19]);
and and372(ip_11_20,x[11],y[20]);
and and373(ip_11_21,x[11],y[21]);
and and374(ip_11_22,x[11],y[22]);
and and375(ip_11_23,x[11],y[23]);
and and376(ip_11_24,x[11],y[24]);
and and377(ip_11_25,x[11],y[25]);
and and378(ip_11_26,x[11],y[26]);
and and379(ip_11_27,x[11],y[27]);
and and380(ip_11_28,x[11],y[28]);
and and381(ip_11_29,x[11],y[29]);
and and382(ip_11_30,x[11],y[30]);
and and383(ip_11_31,x[11],y[31]);
and and384(ip_12_0,x[12],y[0]);
and and385(ip_12_1,x[12],y[1]);
and and386(ip_12_2,x[12],y[2]);
and and387(ip_12_3,x[12],y[3]);
and and388(ip_12_4,x[12],y[4]);
and and389(ip_12_5,x[12],y[5]);
and and390(ip_12_6,x[12],y[6]);
and and391(ip_12_7,x[12],y[7]);
and and392(ip_12_8,x[12],y[8]);
and and393(ip_12_9,x[12],y[9]);
and and394(ip_12_10,x[12],y[10]);
and and395(ip_12_11,x[12],y[11]);
and and396(ip_12_12,x[12],y[12]);
and and397(ip_12_13,x[12],y[13]);
and and398(ip_12_14,x[12],y[14]);
and and399(ip_12_15,x[12],y[15]);
and and400(ip_12_16,x[12],y[16]);
and and401(ip_12_17,x[12],y[17]);
and and402(ip_12_18,x[12],y[18]);
and and403(ip_12_19,x[12],y[19]);
and and404(ip_12_20,x[12],y[20]);
and and405(ip_12_21,x[12],y[21]);
and and406(ip_12_22,x[12],y[22]);
and and407(ip_12_23,x[12],y[23]);
and and408(ip_12_24,x[12],y[24]);
and and409(ip_12_25,x[12],y[25]);
and and410(ip_12_26,x[12],y[26]);
and and411(ip_12_27,x[12],y[27]);
and and412(ip_12_28,x[12],y[28]);
and and413(ip_12_29,x[12],y[29]);
and and414(ip_12_30,x[12],y[30]);
and and415(ip_12_31,x[12],y[31]);
and and416(ip_13_0,x[13],y[0]);
and and417(ip_13_1,x[13],y[1]);
and and418(ip_13_2,x[13],y[2]);
and and419(ip_13_3,x[13],y[3]);
and and420(ip_13_4,x[13],y[4]);
and and421(ip_13_5,x[13],y[5]);
and and422(ip_13_6,x[13],y[6]);
and and423(ip_13_7,x[13],y[7]);
and and424(ip_13_8,x[13],y[8]);
and and425(ip_13_9,x[13],y[9]);
and and426(ip_13_10,x[13],y[10]);
and and427(ip_13_11,x[13],y[11]);
and and428(ip_13_12,x[13],y[12]);
and and429(ip_13_13,x[13],y[13]);
and and430(ip_13_14,x[13],y[14]);
and and431(ip_13_15,x[13],y[15]);
and and432(ip_13_16,x[13],y[16]);
and and433(ip_13_17,x[13],y[17]);
and and434(ip_13_18,x[13],y[18]);
and and435(ip_13_19,x[13],y[19]);
and and436(ip_13_20,x[13],y[20]);
and and437(ip_13_21,x[13],y[21]);
and and438(ip_13_22,x[13],y[22]);
and and439(ip_13_23,x[13],y[23]);
and and440(ip_13_24,x[13],y[24]);
and and441(ip_13_25,x[13],y[25]);
and and442(ip_13_26,x[13],y[26]);
and and443(ip_13_27,x[13],y[27]);
and and444(ip_13_28,x[13],y[28]);
and and445(ip_13_29,x[13],y[29]);
and and446(ip_13_30,x[13],y[30]);
and and447(ip_13_31,x[13],y[31]);
and and448(ip_14_0,x[14],y[0]);
and and449(ip_14_1,x[14],y[1]);
and and450(ip_14_2,x[14],y[2]);
and and451(ip_14_3,x[14],y[3]);
and and452(ip_14_4,x[14],y[4]);
and and453(ip_14_5,x[14],y[5]);
and and454(ip_14_6,x[14],y[6]);
and and455(ip_14_7,x[14],y[7]);
and and456(ip_14_8,x[14],y[8]);
and and457(ip_14_9,x[14],y[9]);
and and458(ip_14_10,x[14],y[10]);
and and459(ip_14_11,x[14],y[11]);
and and460(ip_14_12,x[14],y[12]);
and and461(ip_14_13,x[14],y[13]);
and and462(ip_14_14,x[14],y[14]);
and and463(ip_14_15,x[14],y[15]);
and and464(ip_14_16,x[14],y[16]);
and and465(ip_14_17,x[14],y[17]);
and and466(ip_14_18,x[14],y[18]);
and and467(ip_14_19,x[14],y[19]);
and and468(ip_14_20,x[14],y[20]);
and and469(ip_14_21,x[14],y[21]);
and and470(ip_14_22,x[14],y[22]);
and and471(ip_14_23,x[14],y[23]);
and and472(ip_14_24,x[14],y[24]);
and and473(ip_14_25,x[14],y[25]);
and and474(ip_14_26,x[14],y[26]);
and and475(ip_14_27,x[14],y[27]);
and and476(ip_14_28,x[14],y[28]);
and and477(ip_14_29,x[14],y[29]);
and and478(ip_14_30,x[14],y[30]);
and and479(ip_14_31,x[14],y[31]);
and and480(ip_15_0,x[15],y[0]);
and and481(ip_15_1,x[15],y[1]);
and and482(ip_15_2,x[15],y[2]);
and and483(ip_15_3,x[15],y[3]);
and and484(ip_15_4,x[15],y[4]);
and and485(ip_15_5,x[15],y[5]);
and and486(ip_15_6,x[15],y[6]);
and and487(ip_15_7,x[15],y[7]);
and and488(ip_15_8,x[15],y[8]);
and and489(ip_15_9,x[15],y[9]);
and and490(ip_15_10,x[15],y[10]);
and and491(ip_15_11,x[15],y[11]);
and and492(ip_15_12,x[15],y[12]);
and and493(ip_15_13,x[15],y[13]);
and and494(ip_15_14,x[15],y[14]);
and and495(ip_15_15,x[15],y[15]);
and and496(ip_15_16,x[15],y[16]);
and and497(ip_15_17,x[15],y[17]);
and and498(ip_15_18,x[15],y[18]);
and and499(ip_15_19,x[15],y[19]);
and and500(ip_15_20,x[15],y[20]);
and and501(ip_15_21,x[15],y[21]);
and and502(ip_15_22,x[15],y[22]);
and and503(ip_15_23,x[15],y[23]);
and and504(ip_15_24,x[15],y[24]);
and and505(ip_15_25,x[15],y[25]);
and and506(ip_15_26,x[15],y[26]);
and and507(ip_15_27,x[15],y[27]);
and and508(ip_15_28,x[15],y[28]);
and and509(ip_15_29,x[15],y[29]);
and and510(ip_15_30,x[15],y[30]);
and and511(ip_15_31,x[15],y[31]);
and and512(ip_16_0,x[16],y[0]);
and and513(ip_16_1,x[16],y[1]);
and and514(ip_16_2,x[16],y[2]);
and and515(ip_16_3,x[16],y[3]);
and and516(ip_16_4,x[16],y[4]);
and and517(ip_16_5,x[16],y[5]);
and and518(ip_16_6,x[16],y[6]);
and and519(ip_16_7,x[16],y[7]);
and and520(ip_16_8,x[16],y[8]);
and and521(ip_16_9,x[16],y[9]);
and and522(ip_16_10,x[16],y[10]);
and and523(ip_16_11,x[16],y[11]);
and and524(ip_16_12,x[16],y[12]);
and and525(ip_16_13,x[16],y[13]);
and and526(ip_16_14,x[16],y[14]);
and and527(ip_16_15,x[16],y[15]);
and and528(ip_16_16,x[16],y[16]);
and and529(ip_16_17,x[16],y[17]);
and and530(ip_16_18,x[16],y[18]);
and and531(ip_16_19,x[16],y[19]);
and and532(ip_16_20,x[16],y[20]);
and and533(ip_16_21,x[16],y[21]);
and and534(ip_16_22,x[16],y[22]);
and and535(ip_16_23,x[16],y[23]);
and and536(ip_16_24,x[16],y[24]);
and and537(ip_16_25,x[16],y[25]);
and and538(ip_16_26,x[16],y[26]);
and and539(ip_16_27,x[16],y[27]);
and and540(ip_16_28,x[16],y[28]);
and and541(ip_16_29,x[16],y[29]);
and and542(ip_16_30,x[16],y[30]);
and and543(ip_16_31,x[16],y[31]);
and and544(ip_17_0,x[17],y[0]);
and and545(ip_17_1,x[17],y[1]);
and and546(ip_17_2,x[17],y[2]);
and and547(ip_17_3,x[17],y[3]);
and and548(ip_17_4,x[17],y[4]);
and and549(ip_17_5,x[17],y[5]);
and and550(ip_17_6,x[17],y[6]);
and and551(ip_17_7,x[17],y[7]);
and and552(ip_17_8,x[17],y[8]);
and and553(ip_17_9,x[17],y[9]);
and and554(ip_17_10,x[17],y[10]);
and and555(ip_17_11,x[17],y[11]);
and and556(ip_17_12,x[17],y[12]);
and and557(ip_17_13,x[17],y[13]);
and and558(ip_17_14,x[17],y[14]);
and and559(ip_17_15,x[17],y[15]);
and and560(ip_17_16,x[17],y[16]);
and and561(ip_17_17,x[17],y[17]);
and and562(ip_17_18,x[17],y[18]);
and and563(ip_17_19,x[17],y[19]);
and and564(ip_17_20,x[17],y[20]);
and and565(ip_17_21,x[17],y[21]);
and and566(ip_17_22,x[17],y[22]);
and and567(ip_17_23,x[17],y[23]);
and and568(ip_17_24,x[17],y[24]);
and and569(ip_17_25,x[17],y[25]);
and and570(ip_17_26,x[17],y[26]);
and and571(ip_17_27,x[17],y[27]);
and and572(ip_17_28,x[17],y[28]);
and and573(ip_17_29,x[17],y[29]);
and and574(ip_17_30,x[17],y[30]);
and and575(ip_17_31,x[17],y[31]);
and and576(ip_18_0,x[18],y[0]);
and and577(ip_18_1,x[18],y[1]);
and and578(ip_18_2,x[18],y[2]);
and and579(ip_18_3,x[18],y[3]);
and and580(ip_18_4,x[18],y[4]);
and and581(ip_18_5,x[18],y[5]);
and and582(ip_18_6,x[18],y[6]);
and and583(ip_18_7,x[18],y[7]);
and and584(ip_18_8,x[18],y[8]);
and and585(ip_18_9,x[18],y[9]);
and and586(ip_18_10,x[18],y[10]);
and and587(ip_18_11,x[18],y[11]);
and and588(ip_18_12,x[18],y[12]);
and and589(ip_18_13,x[18],y[13]);
and and590(ip_18_14,x[18],y[14]);
and and591(ip_18_15,x[18],y[15]);
and and592(ip_18_16,x[18],y[16]);
and and593(ip_18_17,x[18],y[17]);
and and594(ip_18_18,x[18],y[18]);
and and595(ip_18_19,x[18],y[19]);
and and596(ip_18_20,x[18],y[20]);
and and597(ip_18_21,x[18],y[21]);
and and598(ip_18_22,x[18],y[22]);
and and599(ip_18_23,x[18],y[23]);
and and600(ip_18_24,x[18],y[24]);
and and601(ip_18_25,x[18],y[25]);
and and602(ip_18_26,x[18],y[26]);
and and603(ip_18_27,x[18],y[27]);
and and604(ip_18_28,x[18],y[28]);
and and605(ip_18_29,x[18],y[29]);
and and606(ip_18_30,x[18],y[30]);
and and607(ip_18_31,x[18],y[31]);
and and608(ip_19_0,x[19],y[0]);
and and609(ip_19_1,x[19],y[1]);
and and610(ip_19_2,x[19],y[2]);
and and611(ip_19_3,x[19],y[3]);
and and612(ip_19_4,x[19],y[4]);
and and613(ip_19_5,x[19],y[5]);
and and614(ip_19_6,x[19],y[6]);
and and615(ip_19_7,x[19],y[7]);
and and616(ip_19_8,x[19],y[8]);
and and617(ip_19_9,x[19],y[9]);
and and618(ip_19_10,x[19],y[10]);
and and619(ip_19_11,x[19],y[11]);
and and620(ip_19_12,x[19],y[12]);
and and621(ip_19_13,x[19],y[13]);
and and622(ip_19_14,x[19],y[14]);
and and623(ip_19_15,x[19],y[15]);
and and624(ip_19_16,x[19],y[16]);
and and625(ip_19_17,x[19],y[17]);
and and626(ip_19_18,x[19],y[18]);
and and627(ip_19_19,x[19],y[19]);
and and628(ip_19_20,x[19],y[20]);
and and629(ip_19_21,x[19],y[21]);
and and630(ip_19_22,x[19],y[22]);
and and631(ip_19_23,x[19],y[23]);
and and632(ip_19_24,x[19],y[24]);
and and633(ip_19_25,x[19],y[25]);
and and634(ip_19_26,x[19],y[26]);
and and635(ip_19_27,x[19],y[27]);
and and636(ip_19_28,x[19],y[28]);
and and637(ip_19_29,x[19],y[29]);
and and638(ip_19_30,x[19],y[30]);
and and639(ip_19_31,x[19],y[31]);
and and640(ip_20_0,x[20],y[0]);
and and641(ip_20_1,x[20],y[1]);
and and642(ip_20_2,x[20],y[2]);
and and643(ip_20_3,x[20],y[3]);
and and644(ip_20_4,x[20],y[4]);
and and645(ip_20_5,x[20],y[5]);
and and646(ip_20_6,x[20],y[6]);
and and647(ip_20_7,x[20],y[7]);
and and648(ip_20_8,x[20],y[8]);
and and649(ip_20_9,x[20],y[9]);
and and650(ip_20_10,x[20],y[10]);
and and651(ip_20_11,x[20],y[11]);
and and652(ip_20_12,x[20],y[12]);
and and653(ip_20_13,x[20],y[13]);
and and654(ip_20_14,x[20],y[14]);
and and655(ip_20_15,x[20],y[15]);
and and656(ip_20_16,x[20],y[16]);
and and657(ip_20_17,x[20],y[17]);
and and658(ip_20_18,x[20],y[18]);
and and659(ip_20_19,x[20],y[19]);
and and660(ip_20_20,x[20],y[20]);
and and661(ip_20_21,x[20],y[21]);
and and662(ip_20_22,x[20],y[22]);
and and663(ip_20_23,x[20],y[23]);
and and664(ip_20_24,x[20],y[24]);
and and665(ip_20_25,x[20],y[25]);
and and666(ip_20_26,x[20],y[26]);
and and667(ip_20_27,x[20],y[27]);
and and668(ip_20_28,x[20],y[28]);
and and669(ip_20_29,x[20],y[29]);
and and670(ip_20_30,x[20],y[30]);
and and671(ip_20_31,x[20],y[31]);
and and672(ip_21_0,x[21],y[0]);
and and673(ip_21_1,x[21],y[1]);
and and674(ip_21_2,x[21],y[2]);
and and675(ip_21_3,x[21],y[3]);
and and676(ip_21_4,x[21],y[4]);
and and677(ip_21_5,x[21],y[5]);
and and678(ip_21_6,x[21],y[6]);
and and679(ip_21_7,x[21],y[7]);
and and680(ip_21_8,x[21],y[8]);
and and681(ip_21_9,x[21],y[9]);
and and682(ip_21_10,x[21],y[10]);
and and683(ip_21_11,x[21],y[11]);
and and684(ip_21_12,x[21],y[12]);
and and685(ip_21_13,x[21],y[13]);
and and686(ip_21_14,x[21],y[14]);
and and687(ip_21_15,x[21],y[15]);
and and688(ip_21_16,x[21],y[16]);
and and689(ip_21_17,x[21],y[17]);
and and690(ip_21_18,x[21],y[18]);
and and691(ip_21_19,x[21],y[19]);
and and692(ip_21_20,x[21],y[20]);
and and693(ip_21_21,x[21],y[21]);
and and694(ip_21_22,x[21],y[22]);
and and695(ip_21_23,x[21],y[23]);
and and696(ip_21_24,x[21],y[24]);
and and697(ip_21_25,x[21],y[25]);
and and698(ip_21_26,x[21],y[26]);
and and699(ip_21_27,x[21],y[27]);
and and700(ip_21_28,x[21],y[28]);
and and701(ip_21_29,x[21],y[29]);
and and702(ip_21_30,x[21],y[30]);
and and703(ip_21_31,x[21],y[31]);
and and704(ip_22_0,x[22],y[0]);
and and705(ip_22_1,x[22],y[1]);
and and706(ip_22_2,x[22],y[2]);
and and707(ip_22_3,x[22],y[3]);
and and708(ip_22_4,x[22],y[4]);
and and709(ip_22_5,x[22],y[5]);
and and710(ip_22_6,x[22],y[6]);
and and711(ip_22_7,x[22],y[7]);
and and712(ip_22_8,x[22],y[8]);
and and713(ip_22_9,x[22],y[9]);
and and714(ip_22_10,x[22],y[10]);
and and715(ip_22_11,x[22],y[11]);
and and716(ip_22_12,x[22],y[12]);
and and717(ip_22_13,x[22],y[13]);
and and718(ip_22_14,x[22],y[14]);
and and719(ip_22_15,x[22],y[15]);
and and720(ip_22_16,x[22],y[16]);
and and721(ip_22_17,x[22],y[17]);
and and722(ip_22_18,x[22],y[18]);
and and723(ip_22_19,x[22],y[19]);
and and724(ip_22_20,x[22],y[20]);
and and725(ip_22_21,x[22],y[21]);
and and726(ip_22_22,x[22],y[22]);
and and727(ip_22_23,x[22],y[23]);
and and728(ip_22_24,x[22],y[24]);
and and729(ip_22_25,x[22],y[25]);
and and730(ip_22_26,x[22],y[26]);
and and731(ip_22_27,x[22],y[27]);
and and732(ip_22_28,x[22],y[28]);
and and733(ip_22_29,x[22],y[29]);
and and734(ip_22_30,x[22],y[30]);
and and735(ip_22_31,x[22],y[31]);
and and736(ip_23_0,x[23],y[0]);
and and737(ip_23_1,x[23],y[1]);
and and738(ip_23_2,x[23],y[2]);
and and739(ip_23_3,x[23],y[3]);
and and740(ip_23_4,x[23],y[4]);
and and741(ip_23_5,x[23],y[5]);
and and742(ip_23_6,x[23],y[6]);
and and743(ip_23_7,x[23],y[7]);
and and744(ip_23_8,x[23],y[8]);
and and745(ip_23_9,x[23],y[9]);
and and746(ip_23_10,x[23],y[10]);
and and747(ip_23_11,x[23],y[11]);
and and748(ip_23_12,x[23],y[12]);
and and749(ip_23_13,x[23],y[13]);
and and750(ip_23_14,x[23],y[14]);
and and751(ip_23_15,x[23],y[15]);
and and752(ip_23_16,x[23],y[16]);
and and753(ip_23_17,x[23],y[17]);
and and754(ip_23_18,x[23],y[18]);
and and755(ip_23_19,x[23],y[19]);
and and756(ip_23_20,x[23],y[20]);
and and757(ip_23_21,x[23],y[21]);
and and758(ip_23_22,x[23],y[22]);
and and759(ip_23_23,x[23],y[23]);
and and760(ip_23_24,x[23],y[24]);
and and761(ip_23_25,x[23],y[25]);
and and762(ip_23_26,x[23],y[26]);
and and763(ip_23_27,x[23],y[27]);
and and764(ip_23_28,x[23],y[28]);
and and765(ip_23_29,x[23],y[29]);
and and766(ip_23_30,x[23],y[30]);
and and767(ip_23_31,x[23],y[31]);
and and768(ip_24_0,x[24],y[0]);
and and769(ip_24_1,x[24],y[1]);
and and770(ip_24_2,x[24],y[2]);
and and771(ip_24_3,x[24],y[3]);
and and772(ip_24_4,x[24],y[4]);
and and773(ip_24_5,x[24],y[5]);
and and774(ip_24_6,x[24],y[6]);
and and775(ip_24_7,x[24],y[7]);
and and776(ip_24_8,x[24],y[8]);
and and777(ip_24_9,x[24],y[9]);
and and778(ip_24_10,x[24],y[10]);
and and779(ip_24_11,x[24],y[11]);
and and780(ip_24_12,x[24],y[12]);
and and781(ip_24_13,x[24],y[13]);
and and782(ip_24_14,x[24],y[14]);
and and783(ip_24_15,x[24],y[15]);
and and784(ip_24_16,x[24],y[16]);
and and785(ip_24_17,x[24],y[17]);
and and786(ip_24_18,x[24],y[18]);
and and787(ip_24_19,x[24],y[19]);
and and788(ip_24_20,x[24],y[20]);
and and789(ip_24_21,x[24],y[21]);
and and790(ip_24_22,x[24],y[22]);
and and791(ip_24_23,x[24],y[23]);
and and792(ip_24_24,x[24],y[24]);
and and793(ip_24_25,x[24],y[25]);
and and794(ip_24_26,x[24],y[26]);
and and795(ip_24_27,x[24],y[27]);
and and796(ip_24_28,x[24],y[28]);
and and797(ip_24_29,x[24],y[29]);
and and798(ip_24_30,x[24],y[30]);
and and799(ip_24_31,x[24],y[31]);
and and800(ip_25_0,x[25],y[0]);
and and801(ip_25_1,x[25],y[1]);
and and802(ip_25_2,x[25],y[2]);
and and803(ip_25_3,x[25],y[3]);
and and804(ip_25_4,x[25],y[4]);
and and805(ip_25_5,x[25],y[5]);
and and806(ip_25_6,x[25],y[6]);
and and807(ip_25_7,x[25],y[7]);
and and808(ip_25_8,x[25],y[8]);
and and809(ip_25_9,x[25],y[9]);
and and810(ip_25_10,x[25],y[10]);
and and811(ip_25_11,x[25],y[11]);
and and812(ip_25_12,x[25],y[12]);
and and813(ip_25_13,x[25],y[13]);
and and814(ip_25_14,x[25],y[14]);
and and815(ip_25_15,x[25],y[15]);
and and816(ip_25_16,x[25],y[16]);
and and817(ip_25_17,x[25],y[17]);
and and818(ip_25_18,x[25],y[18]);
and and819(ip_25_19,x[25],y[19]);
and and820(ip_25_20,x[25],y[20]);
and and821(ip_25_21,x[25],y[21]);
and and822(ip_25_22,x[25],y[22]);
and and823(ip_25_23,x[25],y[23]);
and and824(ip_25_24,x[25],y[24]);
and and825(ip_25_25,x[25],y[25]);
and and826(ip_25_26,x[25],y[26]);
and and827(ip_25_27,x[25],y[27]);
and and828(ip_25_28,x[25],y[28]);
and and829(ip_25_29,x[25],y[29]);
and and830(ip_25_30,x[25],y[30]);
and and831(ip_25_31,x[25],y[31]);
and and832(ip_26_0,x[26],y[0]);
and and833(ip_26_1,x[26],y[1]);
and and834(ip_26_2,x[26],y[2]);
and and835(ip_26_3,x[26],y[3]);
and and836(ip_26_4,x[26],y[4]);
and and837(ip_26_5,x[26],y[5]);
and and838(ip_26_6,x[26],y[6]);
and and839(ip_26_7,x[26],y[7]);
and and840(ip_26_8,x[26],y[8]);
and and841(ip_26_9,x[26],y[9]);
and and842(ip_26_10,x[26],y[10]);
and and843(ip_26_11,x[26],y[11]);
and and844(ip_26_12,x[26],y[12]);
and and845(ip_26_13,x[26],y[13]);
and and846(ip_26_14,x[26],y[14]);
and and847(ip_26_15,x[26],y[15]);
and and848(ip_26_16,x[26],y[16]);
and and849(ip_26_17,x[26],y[17]);
and and850(ip_26_18,x[26],y[18]);
and and851(ip_26_19,x[26],y[19]);
and and852(ip_26_20,x[26],y[20]);
and and853(ip_26_21,x[26],y[21]);
and and854(ip_26_22,x[26],y[22]);
and and855(ip_26_23,x[26],y[23]);
and and856(ip_26_24,x[26],y[24]);
and and857(ip_26_25,x[26],y[25]);
and and858(ip_26_26,x[26],y[26]);
and and859(ip_26_27,x[26],y[27]);
and and860(ip_26_28,x[26],y[28]);
and and861(ip_26_29,x[26],y[29]);
and and862(ip_26_30,x[26],y[30]);
and and863(ip_26_31,x[26],y[31]);
and and864(ip_27_0,x[27],y[0]);
and and865(ip_27_1,x[27],y[1]);
and and866(ip_27_2,x[27],y[2]);
and and867(ip_27_3,x[27],y[3]);
and and868(ip_27_4,x[27],y[4]);
and and869(ip_27_5,x[27],y[5]);
and and870(ip_27_6,x[27],y[6]);
and and871(ip_27_7,x[27],y[7]);
and and872(ip_27_8,x[27],y[8]);
and and873(ip_27_9,x[27],y[9]);
and and874(ip_27_10,x[27],y[10]);
and and875(ip_27_11,x[27],y[11]);
and and876(ip_27_12,x[27],y[12]);
and and877(ip_27_13,x[27],y[13]);
and and878(ip_27_14,x[27],y[14]);
and and879(ip_27_15,x[27],y[15]);
and and880(ip_27_16,x[27],y[16]);
and and881(ip_27_17,x[27],y[17]);
and and882(ip_27_18,x[27],y[18]);
and and883(ip_27_19,x[27],y[19]);
and and884(ip_27_20,x[27],y[20]);
and and885(ip_27_21,x[27],y[21]);
and and886(ip_27_22,x[27],y[22]);
and and887(ip_27_23,x[27],y[23]);
and and888(ip_27_24,x[27],y[24]);
and and889(ip_27_25,x[27],y[25]);
and and890(ip_27_26,x[27],y[26]);
and and891(ip_27_27,x[27],y[27]);
and and892(ip_27_28,x[27],y[28]);
and and893(ip_27_29,x[27],y[29]);
and and894(ip_27_30,x[27],y[30]);
and and895(ip_27_31,x[27],y[31]);
and and896(ip_28_0,x[28],y[0]);
and and897(ip_28_1,x[28],y[1]);
and and898(ip_28_2,x[28],y[2]);
and and899(ip_28_3,x[28],y[3]);
and and900(ip_28_4,x[28],y[4]);
and and901(ip_28_5,x[28],y[5]);
and and902(ip_28_6,x[28],y[6]);
and and903(ip_28_7,x[28],y[7]);
and and904(ip_28_8,x[28],y[8]);
and and905(ip_28_9,x[28],y[9]);
and and906(ip_28_10,x[28],y[10]);
and and907(ip_28_11,x[28],y[11]);
and and908(ip_28_12,x[28],y[12]);
and and909(ip_28_13,x[28],y[13]);
and and910(ip_28_14,x[28],y[14]);
and and911(ip_28_15,x[28],y[15]);
and and912(ip_28_16,x[28],y[16]);
and and913(ip_28_17,x[28],y[17]);
and and914(ip_28_18,x[28],y[18]);
and and915(ip_28_19,x[28],y[19]);
and and916(ip_28_20,x[28],y[20]);
and and917(ip_28_21,x[28],y[21]);
and and918(ip_28_22,x[28],y[22]);
and and919(ip_28_23,x[28],y[23]);
and and920(ip_28_24,x[28],y[24]);
and and921(ip_28_25,x[28],y[25]);
and and922(ip_28_26,x[28],y[26]);
and and923(ip_28_27,x[28],y[27]);
and and924(ip_28_28,x[28],y[28]);
and and925(ip_28_29,x[28],y[29]);
and and926(ip_28_30,x[28],y[30]);
and and927(ip_28_31,x[28],y[31]);
and and928(ip_29_0,x[29],y[0]);
and and929(ip_29_1,x[29],y[1]);
and and930(ip_29_2,x[29],y[2]);
and and931(ip_29_3,x[29],y[3]);
and and932(ip_29_4,x[29],y[4]);
and and933(ip_29_5,x[29],y[5]);
and and934(ip_29_6,x[29],y[6]);
and and935(ip_29_7,x[29],y[7]);
and and936(ip_29_8,x[29],y[8]);
and and937(ip_29_9,x[29],y[9]);
and and938(ip_29_10,x[29],y[10]);
and and939(ip_29_11,x[29],y[11]);
and and940(ip_29_12,x[29],y[12]);
and and941(ip_29_13,x[29],y[13]);
and and942(ip_29_14,x[29],y[14]);
and and943(ip_29_15,x[29],y[15]);
and and944(ip_29_16,x[29],y[16]);
and and945(ip_29_17,x[29],y[17]);
and and946(ip_29_18,x[29],y[18]);
and and947(ip_29_19,x[29],y[19]);
and and948(ip_29_20,x[29],y[20]);
and and949(ip_29_21,x[29],y[21]);
and and950(ip_29_22,x[29],y[22]);
and and951(ip_29_23,x[29],y[23]);
and and952(ip_29_24,x[29],y[24]);
and and953(ip_29_25,x[29],y[25]);
and and954(ip_29_26,x[29],y[26]);
and and955(ip_29_27,x[29],y[27]);
and and956(ip_29_28,x[29],y[28]);
and and957(ip_29_29,x[29],y[29]);
and and958(ip_29_30,x[29],y[30]);
and and959(ip_29_31,x[29],y[31]);
and and960(ip_30_0,x[30],y[0]);
and and961(ip_30_1,x[30],y[1]);
and and962(ip_30_2,x[30],y[2]);
and and963(ip_30_3,x[30],y[3]);
and and964(ip_30_4,x[30],y[4]);
and and965(ip_30_5,x[30],y[5]);
and and966(ip_30_6,x[30],y[6]);
and and967(ip_30_7,x[30],y[7]);
and and968(ip_30_8,x[30],y[8]);
and and969(ip_30_9,x[30],y[9]);
and and970(ip_30_10,x[30],y[10]);
and and971(ip_30_11,x[30],y[11]);
and and972(ip_30_12,x[30],y[12]);
and and973(ip_30_13,x[30],y[13]);
and and974(ip_30_14,x[30],y[14]);
and and975(ip_30_15,x[30],y[15]);
and and976(ip_30_16,x[30],y[16]);
and and977(ip_30_17,x[30],y[17]);
and and978(ip_30_18,x[30],y[18]);
and and979(ip_30_19,x[30],y[19]);
and and980(ip_30_20,x[30],y[20]);
and and981(ip_30_21,x[30],y[21]);
and and982(ip_30_22,x[30],y[22]);
and and983(ip_30_23,x[30],y[23]);
and and984(ip_30_24,x[30],y[24]);
and and985(ip_30_25,x[30],y[25]);
and and986(ip_30_26,x[30],y[26]);
and and987(ip_30_27,x[30],y[27]);
and and988(ip_30_28,x[30],y[28]);
and and989(ip_30_29,x[30],y[29]);
and and990(ip_30_30,x[30],y[30]);
and and991(ip_30_31,x[30],y[31]);
and and992(ip_31_0,x[31],y[0]);
and and993(ip_31_1,x[31],y[1]);
and and994(ip_31_2,x[31],y[2]);
and and995(ip_31_3,x[31],y[3]);
and and996(ip_31_4,x[31],y[4]);
and and997(ip_31_5,x[31],y[5]);
and and998(ip_31_6,x[31],y[6]);
and and999(ip_31_7,x[31],y[7]);
and and1000(ip_31_8,x[31],y[8]);
and and1001(ip_31_9,x[31],y[9]);
and and1002(ip_31_10,x[31],y[10]);
and and1003(ip_31_11,x[31],y[11]);
and and1004(ip_31_12,x[31],y[12]);
and and1005(ip_31_13,x[31],y[13]);
and and1006(ip_31_14,x[31],y[14]);
and and1007(ip_31_15,x[31],y[15]);
and and1008(ip_31_16,x[31],y[16]);
and and1009(ip_31_17,x[31],y[17]);
and and1010(ip_31_18,x[31],y[18]);
and and1011(ip_31_19,x[31],y[19]);
and and1012(ip_31_20,x[31],y[20]);
and and1013(ip_31_21,x[31],y[21]);
and and1014(ip_31_22,x[31],y[22]);
and and1015(ip_31_23,x[31],y[23]);
and and1016(ip_31_24,x[31],y[24]);
and and1017(ip_31_25,x[31],y[25]);
and and1018(ip_31_26,x[31],y[26]);
and and1019(ip_31_27,x[31],y[27]);
and and1020(ip_31_28,x[31],y[28]);
and and1021(ip_31_29,x[31],y[29]);
and and1022(ip_31_30,x[31],y[30]);
and and1023(ip_31_31,x[31],y[31]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
FA fa2(ip_3_0,p3,p0,p4,p5);
FA fa3(ip_0_4,ip_1_3,ip_2_2,p6,p7);
FA fa4(ip_3_1,ip_4_0,p7,p8,p9);
FA fa5(p2,p9,p4,p10,p11);
FA fa6(ip_0_5,ip_1_4,ip_2_3,p12,p13);
FA fa7(ip_3_2,ip_4_1,ip_5_0,p14,p15);
FA fa8(p13,p15,p6,p16,p17);
FA fa9(p17,p8,p10,p18,p19);
FA fa10(ip_0_6,ip_1_5,ip_2_4,p20,p21);
FA fa11(ip_3_3,ip_4_2,ip_5_1,p22,p23);
FA fa12(ip_6_0,p21,p23,p24,p25);
FA fa13(p12,p14,p25,p26,p27);
FA fa14(p16,p27,p18,p28,p29);
FA fa15(ip_0_7,ip_1_6,ip_2_5,p30,p31);
FA fa16(ip_3_4,ip_4_3,ip_5_2,p32,p33);
FA fa17(ip_6_1,ip_7_0,p31,p34,p35);
FA fa18(p33,p20,p22,p36,p37);
FA fa19(p35,p24,p37,p38,p39);
FA fa20(p26,p39,p28,p40,p41);
FA fa21(ip_0_8,ip_1_7,ip_2_6,p42,p43);
FA fa22(ip_3_5,ip_4_4,ip_5_3,p44,p45);
FA fa23(ip_6_2,ip_7_1,ip_8_0,p46,p47);
FA fa24(p43,p45,p47,p48,p49);
FA fa25(p30,p32,p34,p50,p51);
FA fa26(p49,p51,p36,p52,p53);
FA fa27(p53,p38,p40,p54,p55);
FA fa28(ip_0_9,ip_1_8,ip_2_7,p56,p57);
FA fa29(ip_3_6,ip_4_5,ip_5_4,p58,p59);
FA fa30(ip_6_3,ip_7_2,ip_8_1,p60,p61);
FA fa31(ip_9_0,p57,p59,p62,p63);
FA fa32(p61,p42,p44,p64,p65);
FA fa33(p46,p63,p48,p66,p67);
FA fa34(p65,p50,p67,p68,p69);
FA fa35(p52,p69,p54,p70,p71);
FA fa36(ip_0_10,ip_1_9,ip_2_8,p72,p73);
FA fa37(ip_3_7,ip_4_6,ip_5_5,p74,p75);
FA fa38(ip_6_4,ip_7_3,ip_8_2,p76,p77);
FA fa39(ip_9_1,ip_10_0,p73,p78,p79);
FA fa40(p75,p77,p56,p80,p81);
FA fa41(p58,p60,p79,p82,p83);
FA fa42(p81,p62,p83,p84,p85);
FA fa43(p64,p66,p85,p86,p87);
FA fa44(p68,p87,p70,p88,p89);
FA fa45(ip_0_11,ip_1_10,ip_2_9,p90,p91);
FA fa46(ip_3_8,ip_4_7,ip_5_6,p92,p93);
FA fa47(ip_6_5,ip_7_4,ip_8_3,p94,p95);
FA fa48(ip_9_2,ip_10_1,ip_11_0,p96,p97);
FA fa49(p91,p93,p95,p98,p99);
FA fa50(p97,p72,p74,p100,p101);
FA fa51(p76,p78,p99,p102,p103);
FA fa52(p101,p80,p103,p104,p105);
FA fa53(p82,p105,p84,p106,p107);
FA fa54(p107,p86,p88,p108,p109);
FA fa55(ip_0_12,ip_1_11,ip_2_10,p110,p111);
FA fa56(ip_3_9,ip_4_8,ip_5_7,p112,p113);
FA fa57(ip_6_6,ip_7_5,ip_8_4,p114,p115);
FA fa58(ip_9_3,ip_10_2,ip_11_1,p116,p117);
FA fa59(ip_12_0,p111,p113,p118,p119);
FA fa60(p115,p117,p90,p120,p121);
FA fa61(p92,p94,p96,p122,p123);
FA fa62(p119,p121,p123,p124,p125);
FA fa63(p98,p100,p125,p126,p127);
FA fa64(p102,p104,p127,p128,p129);
FA fa65(p106,p129,p108,p130,p131);
FA fa66(ip_0_13,ip_1_12,ip_2_11,p132,p133);
FA fa67(ip_3_10,ip_4_9,ip_5_8,p134,p135);
FA fa68(ip_6_7,ip_7_6,ip_8_5,p136,p137);
FA fa69(ip_9_4,ip_10_3,ip_11_2,p138,p139);
FA fa70(ip_12_1,ip_13_0,p133,p140,p141);
FA fa71(p135,p137,p139,p142,p143);
FA fa72(p110,p112,p114,p144,p145);
FA fa73(p116,p141,p143,p146,p147);
FA fa74(p118,p120,p145,p148,p149);
FA fa75(p147,p122,p124,p150,p151);
FA fa76(p149,p151,p126,p152,p153);
FA fa77(p153,p128,p130,p154,p155);
FA fa78(ip_0_14,ip_1_13,ip_2_12,p156,p157);
FA fa79(ip_3_11,ip_4_10,ip_5_9,p158,p159);
FA fa80(ip_6_8,ip_7_7,ip_8_6,p160,p161);
FA fa81(ip_9_5,ip_10_4,ip_11_3,p162,p163);
FA fa82(ip_12_2,ip_13_1,ip_14_0,p164,p165);
FA fa83(p157,p159,p161,p166,p167);
FA fa84(p163,p165,p132,p168,p169);
FA fa85(p134,p136,p138,p170,p171);
FA fa86(p140,p167,p169,p172,p173);
FA fa87(p142,p171,p144,p174,p175);
FA fa88(p146,p173,p175,p176,p177);
FA fa89(p148,p177,p150,p178,p179);
FA fa90(p179,p152,p154,p180,p181);
FA fa91(ip_0_15,ip_1_14,ip_2_13,p182,p183);
FA fa92(ip_3_12,ip_4_11,ip_5_10,p184,p185);
FA fa93(ip_6_9,ip_7_8,ip_8_7,p186,p187);
FA fa94(ip_9_6,ip_10_5,ip_11_4,p188,p189);
FA fa95(ip_12_3,ip_13_2,ip_14_1,p190,p191);
FA fa96(ip_15_0,p183,p185,p192,p193);
FA fa97(p187,p189,p191,p194,p195);
FA fa98(p156,p158,p160,p196,p197);
FA fa99(p162,p164,p193,p198,p199);
FA fa100(p195,p166,p168,p200,p201);
FA fa101(p197,p199,p170,p202,p203);
FA fa102(p172,p201,p203,p204,p205);
FA fa103(p174,p176,p205,p206,p207);
FA fa104(p178,p207,p180,p208,p209);
FA fa105(ip_0_16,ip_1_15,ip_2_14,p210,p211);
FA fa106(ip_3_13,ip_4_12,ip_5_11,p212,p213);
FA fa107(ip_6_10,ip_7_9,ip_8_8,p214,p215);
FA fa108(ip_9_7,ip_10_6,ip_11_5,p216,p217);
FA fa109(ip_12_4,ip_13_3,ip_14_2,p218,p219);
FA fa110(ip_15_1,ip_16_0,p211,p220,p221);
FA fa111(p213,p215,p217,p222,p223);
FA fa112(p219,p182,p184,p224,p225);
FA fa113(p186,p188,p190,p226,p227);
FA fa114(p221,p223,p192,p228,p229);
FA fa115(p194,p225,p227,p230,p231);
FA fa116(p196,p198,p229,p232,p233);
FA fa117(p231,p200,p202,p234,p235);
FA fa118(p233,p204,p235,p236,p237);
FA fa119(p206,p237,p208,p238,p239);
FA fa120(ip_0_17,ip_1_16,ip_2_15,p240,p241);
FA fa121(ip_3_14,ip_4_13,ip_5_12,p242,p243);
FA fa122(ip_6_11,ip_7_10,ip_8_9,p244,p245);
FA fa123(ip_9_8,ip_10_7,ip_11_6,p246,p247);
FA fa124(ip_12_5,ip_13_4,ip_14_3,p248,p249);
FA fa125(ip_15_2,ip_16_1,ip_17_0,p250,p251);
FA fa126(p241,p243,p245,p252,p253);
FA fa127(p247,p249,p251,p254,p255);
FA fa128(p210,p212,p214,p256,p257);
FA fa129(p216,p218,p220,p258,p259);
FA fa130(p253,p255,p222,p260,p261);
FA fa131(p257,p259,p224,p262,p263);
FA fa132(p226,p261,p228,p264,p265);
FA fa133(p263,p230,p265,p266,p267);
FA fa134(p232,p267,p234,p268,p269);
FA fa135(p269,p236,p238,p270,p271);
FA fa136(ip_0_18,ip_1_17,ip_2_16,p272,p273);
FA fa137(ip_3_15,ip_4_14,ip_5_13,p274,p275);
FA fa138(ip_6_12,ip_7_11,ip_8_10,p276,p277);
FA fa139(ip_9_9,ip_10_8,ip_11_7,p278,p279);
FA fa140(ip_12_6,ip_13_5,ip_14_4,p280,p281);
FA fa141(ip_15_3,ip_16_2,ip_17_1,p282,p283);
FA fa142(ip_18_0,p273,p275,p284,p285);
FA fa143(p277,p279,p281,p286,p287);
FA fa144(p283,p240,p242,p288,p289);
FA fa145(p244,p246,p248,p290,p291);
FA fa146(p250,p285,p287,p292,p293);
FA fa147(p252,p254,p289,p294,p295);
FA fa148(p291,p256,p258,p296,p297);
FA fa149(p293,p260,p295,p298,p299);
FA fa150(p262,p297,p264,p300,p301);
FA fa151(p299,p301,p266,p302,p303);
FA fa152(p303,p268,p270,p304,p305);
FA fa153(ip_0_19,ip_1_18,ip_2_17,p306,p307);
FA fa154(ip_3_16,ip_4_15,ip_5_14,p308,p309);
FA fa155(ip_6_13,ip_7_12,ip_8_11,p310,p311);
FA fa156(ip_9_10,ip_10_9,ip_11_8,p312,p313);
FA fa157(ip_12_7,ip_13_6,ip_14_5,p314,p315);
FA fa158(ip_15_4,ip_16_3,ip_17_2,p316,p317);
FA fa159(ip_18_1,ip_19_0,p307,p318,p319);
FA fa160(p309,p311,p313,p320,p321);
FA fa161(p315,p317,p272,p322,p323);
FA fa162(p274,p276,p278,p324,p325);
FA fa163(p280,p282,p319,p326,p327);
FA fa164(p321,p323,p284,p328,p329);
FA fa165(p286,p325,p327,p330,p331);
FA fa166(p288,p290,p329,p332,p333);
FA fa167(p292,p331,p294,p334,p335);
FA fa168(p333,p296,p335,p336,p337);
FA fa169(p298,p300,p337,p338,p339);
FA fa170(p302,p339,p304,p340,p341);
FA fa171(ip_0_20,ip_1_19,ip_2_18,p342,p343);
FA fa172(ip_3_17,ip_4_16,ip_5_15,p344,p345);
FA fa173(ip_6_14,ip_7_13,ip_8_12,p346,p347);
FA fa174(ip_9_11,ip_10_10,ip_11_9,p348,p349);
FA fa175(ip_12_8,ip_13_7,ip_14_6,p350,p351);
FA fa176(ip_15_5,ip_16_4,ip_17_3,p352,p353);
FA fa177(ip_18_2,ip_19_1,ip_20_0,p354,p355);
FA fa178(p343,p345,p347,p356,p357);
FA fa179(p349,p351,p353,p358,p359);
FA fa180(p355,p306,p308,p360,p361);
FA fa181(p310,p312,p314,p362,p363);
FA fa182(p316,p318,p357,p364,p365);
FA fa183(p359,p320,p322,p366,p367);
FA fa184(p361,p363,p324,p368,p369);
FA fa185(p326,p365,p328,p370,p371);
FA fa186(p367,p369,p330,p372,p373);
FA fa187(p371,p332,p373,p374,p375);
FA fa188(p334,p375,p336,p376,p377);
FA fa189(p377,p338,p340,p378,p379);
FA fa190(ip_0_21,ip_1_20,ip_2_19,p380,p381);
FA fa191(ip_3_18,ip_4_17,ip_5_16,p382,p383);
FA fa192(ip_6_15,ip_7_14,ip_8_13,p384,p385);
FA fa193(ip_9_12,ip_10_11,ip_11_10,p386,p387);
FA fa194(ip_12_9,ip_13_8,ip_14_7,p388,p389);
FA fa195(ip_15_6,ip_16_5,ip_17_4,p390,p391);
FA fa196(ip_18_3,ip_19_2,ip_20_1,p392,p393);
FA fa197(ip_21_0,p381,p383,p394,p395);
FA fa198(p385,p387,p389,p396,p397);
FA fa199(p391,p393,p342,p398,p399);
FA fa200(p344,p346,p348,p400,p401);
FA fa201(p350,p352,p354,p402,p403);
FA fa202(p395,p397,p399,p404,p405);
FA fa203(p356,p358,p401,p406,p407);
FA fa204(p403,p360,p362,p408,p409);
FA fa205(p405,p364,p407,p410,p411);
FA fa206(p366,p368,p409,p412,p413);
FA fa207(p370,p411,p372,p414,p415);
FA fa208(p413,p415,p374,p416,p417);
FA fa209(p417,p376,p378,p418,p419);
FA fa210(ip_0_22,ip_1_21,ip_2_20,p420,p421);
FA fa211(ip_3_19,ip_4_18,ip_5_17,p422,p423);
FA fa212(ip_6_16,ip_7_15,ip_8_14,p424,p425);
FA fa213(ip_9_13,ip_10_12,ip_11_11,p426,p427);
FA fa214(ip_12_10,ip_13_9,ip_14_8,p428,p429);
FA fa215(ip_15_7,ip_16_6,ip_17_5,p430,p431);
FA fa216(ip_18_4,ip_19_3,ip_20_2,p432,p433);
FA fa217(ip_21_1,ip_22_0,p421,p434,p435);
FA fa218(p423,p425,p427,p436,p437);
FA fa219(p429,p431,p433,p438,p439);
FA fa220(p380,p382,p384,p440,p441);
FA fa221(p386,p388,p390,p442,p443);
FA fa222(p392,p435,p437,p444,p445);
FA fa223(p439,p394,p396,p446,p447);
FA fa224(p398,p441,p443,p448,p449);
FA fa225(p445,p400,p402,p450,p451);
FA fa226(p404,p447,p449,p452,p453);
FA fa227(p406,p451,p408,p454,p455);
FA fa228(p453,p410,p455,p456,p457);
FA fa229(p412,p414,p457,p458,p459);
FA fa230(p416,p459,p418,p460,p461);
FA fa231(ip_0_23,ip_1_22,ip_2_21,p462,p463);
FA fa232(ip_3_20,ip_4_19,ip_5_18,p464,p465);
FA fa233(ip_6_17,ip_7_16,ip_8_15,p466,p467);
FA fa234(ip_9_14,ip_10_13,ip_11_12,p468,p469);
FA fa235(ip_12_11,ip_13_10,ip_14_9,p470,p471);
FA fa236(ip_15_8,ip_16_7,ip_17_6,p472,p473);
FA fa237(ip_18_5,ip_19_4,ip_20_3,p474,p475);
FA fa238(ip_21_2,ip_22_1,ip_23_0,p476,p477);
FA fa239(p463,p465,p467,p478,p479);
FA fa240(p469,p471,p473,p480,p481);
FA fa241(p475,p477,p420,p482,p483);
FA fa242(p422,p424,p426,p484,p485);
FA fa243(p428,p430,p432,p486,p487);
FA fa244(p434,p479,p481,p488,p489);
FA fa245(p483,p436,p438,p490,p491);
FA fa246(p485,p487,p440,p492,p493);
FA fa247(p442,p444,p489,p494,p495);
FA fa248(p491,p493,p446,p496,p497);
FA fa249(p448,p495,p450,p498,p499);
FA fa250(p497,p452,p499,p500,p501);
FA fa251(p454,p501,p456,p502,p503);
FA fa252(p503,p458,p460,p504,p505);
FA fa253(ip_0_24,ip_1_23,ip_2_22,p506,p507);
FA fa254(ip_3_21,ip_4_20,ip_5_19,p508,p509);
FA fa255(ip_6_18,ip_7_17,ip_8_16,p510,p511);
FA fa256(ip_9_15,ip_10_14,ip_11_13,p512,p513);
FA fa257(ip_12_12,ip_13_11,ip_14_10,p514,p515);
FA fa258(ip_15_9,ip_16_8,ip_17_7,p516,p517);
FA fa259(ip_18_6,ip_19_5,ip_20_4,p518,p519);
FA fa260(ip_21_3,ip_22_2,ip_23_1,p520,p521);
FA fa261(ip_24_0,p507,p509,p522,p523);
FA fa262(p511,p513,p515,p524,p525);
FA fa263(p517,p519,p521,p526,p527);
FA fa264(p462,p464,p466,p528,p529);
FA fa265(p468,p470,p472,p530,p531);
FA fa266(p474,p476,p523,p532,p533);
FA fa267(p525,p527,p478,p534,p535);
FA fa268(p480,p482,p529,p536,p537);
FA fa269(p531,p533,p484,p538,p539);
FA fa270(p486,p535,p488,p540,p541);
FA fa271(p537,p539,p490,p542,p543);
FA fa272(p492,p541,p494,p544,p545);
FA fa273(p543,p496,p545,p546,p547);
FA fa274(p498,p547,p500,p548,p549);
FA fa275(p549,p502,p504,p550,p551);
FA fa276(ip_0_25,ip_1_24,ip_2_23,p552,p553);
FA fa277(ip_3_22,ip_4_21,ip_5_20,p554,p555);
FA fa278(ip_6_19,ip_7_18,ip_8_17,p556,p557);
FA fa279(ip_9_16,ip_10_15,ip_11_14,p558,p559);
FA fa280(ip_12_13,ip_13_12,ip_14_11,p560,p561);
FA fa281(ip_15_10,ip_16_9,ip_17_8,p562,p563);
FA fa282(ip_18_7,ip_19_6,ip_20_5,p564,p565);
FA fa283(ip_21_4,ip_22_3,ip_23_2,p566,p567);
FA fa284(ip_24_1,ip_25_0,p553,p568,p569);
FA fa285(p555,p557,p559,p570,p571);
FA fa286(p561,p563,p565,p572,p573);
FA fa287(p567,p506,p508,p574,p575);
FA fa288(p510,p512,p514,p576,p577);
FA fa289(p516,p518,p520,p578,p579);
FA fa290(p569,p571,p573,p580,p581);
FA fa291(p522,p524,p526,p582,p583);
FA fa292(p575,p577,p579,p584,p585);
FA fa293(p528,p530,p532,p586,p587);
FA fa294(p581,p534,p583,p588,p589);
FA fa295(p585,p536,p538,p590,p591);
FA fa296(p587,p540,p589,p592,p593);
FA fa297(p542,p591,p544,p594,p595);
FA fa298(p593,p595,p546,p596,p597);
FA fa299(p597,p548,p550,p598,p599);
FA fa300(ip_0_26,ip_1_25,ip_2_24,p600,p601);
FA fa301(ip_3_23,ip_4_22,ip_5_21,p602,p603);
FA fa302(ip_6_20,ip_7_19,ip_8_18,p604,p605);
FA fa303(ip_9_17,ip_10_16,ip_11_15,p606,p607);
FA fa304(ip_12_14,ip_13_13,ip_14_12,p608,p609);
FA fa305(ip_15_11,ip_16_10,ip_17_9,p610,p611);
FA fa306(ip_18_8,ip_19_7,ip_20_6,p612,p613);
FA fa307(ip_21_5,ip_22_4,ip_23_3,p614,p615);
FA fa308(ip_24_2,ip_25_1,ip_26_0,p616,p617);
FA fa309(p601,p603,p605,p618,p619);
FA fa310(p607,p609,p611,p620,p621);
FA fa311(p613,p615,p617,p622,p623);
FA fa312(p552,p554,p556,p624,p625);
FA fa313(p558,p560,p562,p626,p627);
FA fa314(p564,p566,p568,p628,p629);
FA fa315(p619,p621,p623,p630,p631);
FA fa316(p570,p572,p625,p632,p633);
FA fa317(p627,p629,p574,p634,p635);
FA fa318(p576,p578,p631,p636,p637);
FA fa319(p580,p633,p635,p638,p639);
FA fa320(p582,p584,p637,p640,p641);
FA fa321(p586,p639,p588,p642,p643);
FA fa322(p641,p590,p643,p644,p645);
FA fa323(p592,p594,p645,p646,p647);
FA fa324(p596,p647,p598,p648,p649);
FA fa325(ip_0_27,ip_1_26,ip_2_25,p650,p651);
FA fa326(ip_3_24,ip_4_23,ip_5_22,p652,p653);
FA fa327(ip_6_21,ip_7_20,ip_8_19,p654,p655);
FA fa328(ip_9_18,ip_10_17,ip_11_16,p656,p657);
FA fa329(ip_12_15,ip_13_14,ip_14_13,p658,p659);
FA fa330(ip_15_12,ip_16_11,ip_17_10,p660,p661);
FA fa331(ip_18_9,ip_19_8,ip_20_7,p662,p663);
FA fa332(ip_21_6,ip_22_5,ip_23_4,p664,p665);
FA fa333(ip_24_3,ip_25_2,ip_26_1,p666,p667);
FA fa334(ip_27_0,p651,p653,p668,p669);
FA fa335(p655,p657,p659,p670,p671);
FA fa336(p661,p663,p665,p672,p673);
FA fa337(p667,p600,p602,p674,p675);
FA fa338(p604,p606,p608,p676,p677);
FA fa339(p610,p612,p614,p678,p679);
FA fa340(p616,p669,p671,p680,p681);
FA fa341(p673,p618,p620,p682,p683);
FA fa342(p622,p675,p677,p684,p685);
FA fa343(p679,p624,p626,p686,p687);
FA fa344(p628,p681,p630,p688,p689);
FA fa345(p683,p685,p632,p690,p691);
FA fa346(p634,p687,p689,p692,p693);
FA fa347(p636,p691,p638,p694,p695);
FA fa348(p693,p640,p695,p696,p697);
FA fa349(p642,p697,p644,p698,p699);
FA fa350(p699,p646,p648,p700,p701);
FA fa351(ip_0_28,ip_1_27,ip_2_26,p702,p703);
FA fa352(ip_3_25,ip_4_24,ip_5_23,p704,p705);
FA fa353(ip_6_22,ip_7_21,ip_8_20,p706,p707);
FA fa354(ip_9_19,ip_10_18,ip_11_17,p708,p709);
FA fa355(ip_12_16,ip_13_15,ip_14_14,p710,p711);
FA fa356(ip_15_13,ip_16_12,ip_17_11,p712,p713);
FA fa357(ip_18_10,ip_19_9,ip_20_8,p714,p715);
FA fa358(ip_21_7,ip_22_6,ip_23_5,p716,p717);
FA fa359(ip_24_4,ip_25_3,ip_26_2,p718,p719);
FA fa360(ip_27_1,ip_28_0,p703,p720,p721);
FA fa361(p705,p707,p709,p722,p723);
FA fa362(p711,p713,p715,p724,p725);
FA fa363(p717,p719,p650,p726,p727);
FA fa364(p652,p654,p656,p728,p729);
FA fa365(p658,p660,p662,p730,p731);
FA fa366(p664,p666,p721,p732,p733);
FA fa367(p723,p725,p727,p734,p735);
FA fa368(p668,p670,p672,p736,p737);
FA fa369(p729,p731,p733,p738,p739);
FA fa370(p674,p676,p678,p740,p741);
FA fa371(p735,p680,p737,p742,p743);
FA fa372(p739,p682,p684,p744,p745);
FA fa373(p741,p686,p688,p746,p747);
FA fa374(p743,p690,p745,p748,p749);
FA fa375(p692,p747,p694,p750,p751);
FA fa376(p749,p751,p696,p752,p753);
FA fa377(p753,p698,p700,p754,p755);
FA fa378(ip_0_29,ip_1_28,ip_2_27,p756,p757);
FA fa379(ip_3_26,ip_4_25,ip_5_24,p758,p759);
FA fa380(ip_6_23,ip_7_22,ip_8_21,p760,p761);
FA fa381(ip_9_20,ip_10_19,ip_11_18,p762,p763);
FA fa382(ip_12_17,ip_13_16,ip_14_15,p764,p765);
FA fa383(ip_15_14,ip_16_13,ip_17_12,p766,p767);
FA fa384(ip_18_11,ip_19_10,ip_20_9,p768,p769);
FA fa385(ip_21_8,ip_22_7,ip_23_6,p770,p771);
FA fa386(ip_24_5,ip_25_4,ip_26_3,p772,p773);
FA fa387(ip_27_2,ip_28_1,ip_29_0,p774,p775);
FA fa388(p757,p759,p761,p776,p777);
FA fa389(p763,p765,p767,p778,p779);
FA fa390(p769,p771,p773,p780,p781);
FA fa391(p775,p702,p704,p782,p783);
FA fa392(p706,p708,p710,p784,p785);
FA fa393(p712,p714,p716,p786,p787);
FA fa394(p718,p720,p777,p788,p789);
FA fa395(p779,p781,p722,p790,p791);
FA fa396(p724,p726,p783,p792,p793);
FA fa397(p785,p787,p728,p794,p795);
HA ha0(p730,p732,p796,p797);
FA fa398(p789,p791,p734,p798,p799);
FA fa399(p793,p795,p797,p800,p801);
FA fa400(p736,p738,p799,p802,p803);
FA fa401(p740,p801,p742,p804,p805);
FA fa402(p803,p744,p805,p806,p807);
FA fa403(p746,p748,p807,p808,p809);
FA fa404(p750,p809,p752,p810,p811);
FA fa405(ip_0_30,ip_1_29,ip_2_28,p812,p813);
FA fa406(ip_3_27,ip_4_26,ip_5_25,p814,p815);
FA fa407(ip_6_24,ip_7_23,ip_8_22,p816,p817);
FA fa408(ip_9_21,ip_10_20,ip_11_19,p818,p819);
FA fa409(ip_12_18,ip_13_17,ip_14_16,p820,p821);
FA fa410(ip_15_15,ip_16_14,ip_17_13,p822,p823);
FA fa411(ip_18_12,ip_19_11,ip_20_10,p824,p825);
FA fa412(ip_21_9,ip_22_8,ip_23_7,p826,p827);
FA fa413(ip_24_6,ip_25_5,ip_26_4,p828,p829);
FA fa414(ip_27_3,ip_28_2,ip_29_1,p830,p831);
FA fa415(ip_30_0,p813,p815,p832,p833);
FA fa416(p817,p819,p821,p834,p835);
FA fa417(p823,p825,p827,p836,p837);
FA fa418(p829,p831,p756,p838,p839);
FA fa419(p758,p760,p762,p840,p841);
FA fa420(p764,p766,p768,p842,p843);
FA fa421(p770,p772,p774,p844,p845);
FA fa422(p833,p835,p837,p846,p847);
FA fa423(p839,p776,p778,p848,p849);
FA fa424(p780,p841,p843,p850,p851);
FA fa425(p845,p782,p784,p852,p853);
FA fa426(p786,p847,p788,p854,p855);
FA fa427(p790,p796,p849,p856,p857);
FA fa428(p851,p792,p794,p858,p859);
FA fa429(p853,p855,p798,p860,p861);
FA fa430(p857,p800,p859,p862,p863);
FA fa431(p861,p802,p804,p864,p865);
FA fa432(p863,p865,p806,p866,p867);
FA fa433(p867,p808,p810,p868,p869);
FA fa434(ip_0_31,ip_1_30,ip_2_29,p870,p871);
FA fa435(ip_3_28,ip_4_27,ip_5_26,p872,p873);
FA fa436(ip_6_25,ip_7_24,ip_8_23,p874,p875);
FA fa437(ip_9_22,ip_10_21,ip_11_20,p876,p877);
FA fa438(ip_12_19,ip_13_18,ip_14_17,p878,p879);
FA fa439(ip_15_16,ip_16_15,ip_17_14,p880,p881);
FA fa440(ip_18_13,ip_19_12,ip_20_11,p882,p883);
FA fa441(ip_21_10,ip_22_9,ip_23_8,p884,p885);
FA fa442(ip_24_7,ip_25_6,ip_26_5,p886,p887);
FA fa443(ip_27_4,ip_28_3,ip_29_2,p888,p889);
FA fa444(ip_30_1,ip_31_0,p871,p890,p891);
FA fa445(p873,p875,p877,p892,p893);
FA fa446(p879,p881,p883,p894,p895);
FA fa447(p885,p887,p889,p896,p897);
FA fa448(p812,p814,p816,p898,p899);
FA fa449(p818,p820,p822,p900,p901);
FA fa450(p824,p826,p828,p902,p903);
FA fa451(p830,p891,p893,p904,p905);
FA fa452(p895,p897,p832,p906,p907);
FA fa453(p834,p836,p838,p908,p909);
FA fa454(p899,p901,p903,p910,p911);
FA fa455(p905,p840,p842,p912,p913);
FA fa456(p844,p907,p846,p914,p915);
FA fa457(p909,p911,p848,p916,p917);
FA fa458(p850,p913,p915,p918,p919);
FA fa459(p852,p854,p917,p920,p921);
FA fa460(p856,p919,p858,p922,p923);
FA fa461(p860,p921,p923,p924,p925);
FA fa462(p862,p925,p864,p926,p927);
FA fa463(p927,p866,p868,p928,p929);
FA fa464(ip_1_31,ip_2_30,ip_3_29,p930,p931);
FA fa465(ip_4_28,ip_5_27,ip_6_26,p932,p933);
FA fa466(ip_7_25,ip_8_24,ip_9_23,p934,p935);
FA fa467(ip_10_22,ip_11_21,ip_12_20,p936,p937);
FA fa468(ip_13_19,ip_14_18,ip_15_17,p938,p939);
FA fa469(ip_16_16,ip_17_15,ip_18_14,p940,p941);
FA fa470(ip_19_13,ip_20_12,ip_21_11,p942,p943);
FA fa471(ip_22_10,ip_23_9,ip_24_8,p944,p945);
FA fa472(ip_25_7,ip_26_6,ip_27_5,p946,p947);
FA fa473(ip_28_4,ip_29_3,ip_30_2,p948,p949);
FA fa474(ip_31_1,p931,p933,p950,p951);
FA fa475(p935,p937,p939,p952,p953);
FA fa476(p941,p943,p945,p954,p955);
FA fa477(p947,p949,p870,p956,p957);
FA fa478(p872,p874,p876,p958,p959);
FA fa479(p878,p880,p882,p960,p961);
FA fa480(p884,p886,p888,p962,p963);
FA fa481(p890,p951,p953,p964,p965);
FA fa482(p955,p957,p892,p966,p967);
FA fa483(p894,p896,p959,p968,p969);
FA fa484(p961,p963,p898,p970,p971);
FA fa485(p900,p902,p904,p972,p973);
FA fa486(p965,p967,p906,p974,p975);
FA fa487(p969,p971,p908,p976,p977);
FA fa488(p910,p973,p975,p978,p979);
FA fa489(p912,p914,p977,p980,p981);
FA fa490(p916,p979,p918,p982,p983);
FA fa491(p981,p920,p983,p984,p985);
FA fa492(p922,p924,p985,p986,p987);
FA fa493(p926,p987,p928,p988,p989);
FA fa494(ip_2_31,ip_3_30,ip_4_29,p990,p991);
FA fa495(ip_5_28,ip_6_27,ip_7_26,p992,p993);
FA fa496(ip_8_25,ip_9_24,ip_10_23,p994,p995);
FA fa497(ip_11_22,ip_12_21,ip_13_20,p996,p997);
FA fa498(ip_14_19,ip_15_18,ip_16_17,p998,p999);
FA fa499(ip_17_16,ip_18_15,ip_19_14,p1000,p1001);
FA fa500(ip_20_13,ip_21_12,ip_22_11,p1002,p1003);
FA fa501(ip_23_10,ip_24_9,ip_25_8,p1004,p1005);
FA fa502(ip_26_7,ip_27_6,ip_28_5,p1006,p1007);
FA fa503(ip_29_4,ip_30_3,ip_31_2,p1008,p1009);
FA fa504(p1001,p1003,p1005,p1010,p1011);
FA fa505(p1007,p1009,p991,p1012,p1013);
HA ha1(p993,p995,p1014,p1015);
FA fa506(p997,p999,p1015,p1016,p1017);
FA fa507(p930,p932,p934,p1018,p1019);
FA fa508(p936,p938,p940,p1020,p1021);
FA fa509(p942,p944,p946,p1022,p1023);
FA fa510(p948,p1011,p1013,p1024,p1025);
FA fa511(p1017,p1019,p1021,p1026,p1027);
FA fa512(p1023,p950,p952,p1028,p1029);
FA fa513(p954,p956,p1025,p1030,p1031);
FA fa514(p958,p960,p962,p1032,p1033);
FA fa515(p1027,p1029,p1031,p1034,p1035);
FA fa516(p964,p966,p1033,p1036,p1037);
FA fa517(p968,p970,p1035,p1038,p1039);
FA fa518(p1037,p972,p974,p1040,p1041);
FA fa519(p1039,p976,p1041,p1042,p1043);
FA fa520(p978,p1043,p980,p1044,p1045);
FA fa521(p982,p1045,p984,p1046,p1047);
FA fa522(p1047,p986,p988,p1048,p1049);
FA fa523(ip_3_31,ip_4_30,ip_5_29,p1050,p1051);
FA fa524(ip_6_28,ip_7_27,ip_8_26,p1052,p1053);
FA fa525(ip_9_25,ip_10_24,ip_11_23,p1054,p1055);
FA fa526(ip_12_22,ip_13_21,ip_14_20,p1056,p1057);
FA fa527(ip_15_19,ip_16_18,ip_17_17,p1058,p1059);
FA fa528(ip_18_16,ip_19_15,ip_20_14,p1060,p1061);
FA fa529(ip_21_13,ip_22_12,ip_23_11,p1062,p1063);
FA fa530(ip_24_10,ip_25_9,ip_26_8,p1064,p1065);
FA fa531(ip_27_7,ip_28_6,ip_29_5,p1066,p1067);
FA fa532(ip_30_4,ip_31_3,p1051,p1068,p1069);
FA fa533(p1053,p1055,p1057,p1070,p1071);
FA fa534(p1059,p1061,p1063,p1072,p1073);
FA fa535(p1065,p1067,p1000,p1074,p1075);
FA fa536(p1002,p1004,p1006,p1076,p1077);
FA fa537(p1008,p1014,p1069,p1078,p1079);
FA fa538(p990,p992,p994,p1080,p1081);
FA fa539(p996,p998,p1071,p1082,p1083);
FA fa540(p1073,p1075,p1010,p1084,p1085);
FA fa541(p1012,p1016,p1077,p1086,p1087);
FA fa542(p1079,p1081,p1083,p1088,p1089);
FA fa543(p1018,p1020,p1022,p1090,p1091);
FA fa544(p1085,p1024,p1087,p1092,p1093);
FA fa545(p1089,p1026,p1028,p1094,p1095);
FA fa546(p1030,p1091,p1032,p1096,p1097);
FA fa547(p1093,p1034,p1036,p1098,p1099);
FA fa548(p1095,p1097,p1038,p1100,p1101);
FA fa549(p1040,p1099,p1101,p1102,p1103);
FA fa550(p1042,p1103,p1044,p1104,p1105);
FA fa551(p1105,p1046,p1048,p1106,p1107);
FA fa552(ip_4_31,ip_5_30,ip_6_29,p1108,p1109);
FA fa553(ip_7_28,ip_8_27,ip_9_26,p1110,p1111);
FA fa554(ip_10_25,ip_11_24,ip_12_23,p1112,p1113);
FA fa555(ip_13_22,ip_14_21,ip_15_20,p1114,p1115);
FA fa556(ip_16_19,ip_17_18,ip_18_17,p1116,p1117);
FA fa557(ip_19_16,ip_20_15,ip_21_14,p1118,p1119);
FA fa558(ip_22_13,ip_23_12,ip_24_11,p1120,p1121);
FA fa559(ip_25_10,ip_26_9,ip_27_8,p1122,p1123);
FA fa560(ip_28_7,ip_29_6,ip_30_5,p1124,p1125);
FA fa561(ip_31_4,p1109,p1111,p1126,p1127);
FA fa562(p1113,p1115,p1117,p1128,p1129);
FA fa563(p1119,p1121,p1123,p1130,p1131);
FA fa564(p1125,p1050,p1052,p1132,p1133);
FA fa565(p1054,p1056,p1058,p1134,p1135);
FA fa566(p1060,p1062,p1064,p1136,p1137);
FA fa567(p1066,p1068,p1127,p1138,p1139);
FA fa568(p1129,p1131,p1070,p1140,p1141);
FA fa569(p1072,p1074,p1133,p1142,p1143);
FA fa570(p1135,p1137,p1076,p1144,p1145);
FA fa571(p1078,p1080,p1082,p1146,p1147);
FA fa572(p1139,p1141,p1084,p1148,p1149);
FA fa573(p1143,p1145,p1086,p1150,p1151);
FA fa574(p1088,p1147,p1149,p1152,p1153);
FA fa575(p1090,p1151,p1092,p1154,p1155);
FA fa576(p1153,p1094,p1096,p1156,p1157);
FA fa577(p1155,p1098,p1100,p1158,p1159);
FA fa578(p1157,p1102,p1159,p1160,p1161);
FA fa579(p1104,p1161,p1106,p1162,p1163);
FA fa580(ip_5_31,ip_6_30,ip_7_29,p1164,p1165);
FA fa581(ip_8_28,ip_9_27,ip_10_26,p1166,p1167);
FA fa582(ip_11_25,ip_12_24,ip_13_23,p1168,p1169);
FA fa583(ip_14_22,ip_15_21,ip_16_20,p1170,p1171);
FA fa584(ip_17_19,ip_18_18,ip_19_17,p1172,p1173);
FA fa585(ip_20_16,ip_21_15,ip_22_14,p1174,p1175);
FA fa586(ip_23_13,ip_24_12,ip_25_11,p1176,p1177);
FA fa587(ip_26_10,ip_27_9,ip_28_8,p1178,p1179);
FA fa588(ip_29_7,ip_30_6,ip_31_5,p1180,p1181);
FA fa589(p1165,p1167,p1169,p1182,p1183);
FA fa590(p1171,p1173,p1175,p1184,p1185);
FA fa591(p1177,p1179,p1181,p1186,p1187);
FA fa592(p1108,p1110,p1112,p1188,p1189);
FA fa593(p1114,p1116,p1118,p1190,p1191);
FA fa594(p1120,p1122,p1124,p1192,p1193);
FA fa595(p1183,p1185,p1187,p1194,p1195);
FA fa596(p1126,p1128,p1130,p1196,p1197);
FA fa597(p1189,p1191,p1193,p1198,p1199);
FA fa598(p1132,p1134,p1136,p1200,p1201);
FA fa599(p1195,p1138,p1140,p1202,p1203);
FA fa600(p1197,p1199,p1142,p1204,p1205);
FA fa601(p1144,p1201,p1146,p1206,p1207);
FA fa602(p1148,p1203,p1205,p1208,p1209);
FA fa603(p1150,p1207,p1152,p1210,p1211);
FA fa604(p1209,p1154,p1211,p1212,p1213);
FA fa605(p1156,p1213,p1158,p1214,p1215);
FA fa606(p1215,p1160,p1162,p1216,p1217);
FA fa607(ip_6_31,ip_7_30,ip_8_29,p1218,p1219);
FA fa608(ip_9_28,ip_10_27,ip_11_26,p1220,p1221);
FA fa609(ip_12_25,ip_13_24,ip_14_23,p1222,p1223);
FA fa610(ip_15_22,ip_16_21,ip_17_20,p1224,p1225);
FA fa611(ip_18_19,ip_19_18,ip_20_17,p1226,p1227);
FA fa612(ip_21_16,ip_22_15,ip_23_14,p1228,p1229);
FA fa613(ip_24_13,ip_25_12,ip_26_11,p1230,p1231);
FA fa614(ip_27_10,ip_28_9,ip_29_8,p1232,p1233);
FA fa615(ip_30_7,ip_31_6,p1219,p1234,p1235);
FA fa616(p1221,p1223,p1225,p1236,p1237);
FA fa617(p1227,p1229,p1231,p1238,p1239);
FA fa618(p1233,p1164,p1166,p1240,p1241);
FA fa619(p1168,p1170,p1172,p1242,p1243);
FA fa620(p1174,p1176,p1178,p1244,p1245);
FA fa621(p1180,p1235,p1237,p1246,p1247);
FA fa622(p1239,p1182,p1184,p1248,p1249);
FA fa623(p1186,p1241,p1243,p1250,p1251);
FA fa624(p1245,p1247,p1188,p1252,p1253);
FA fa625(p1190,p1192,p1194,p1254,p1255);
FA fa626(p1249,p1251,p1253,p1256,p1257);
FA fa627(p1196,p1198,p1255,p1258,p1259);
FA fa628(p1200,p1257,p1202,p1260,p1261);
FA fa629(p1204,p1259,p1206,p1262,p1263);
FA fa630(p1261,p1208,p1263,p1264,p1265);
FA fa631(p1210,p1265,p1212,p1266,p1267);
FA fa632(p1267,p1214,p1216,p1268,p1269);
FA fa633(ip_7_31,ip_8_30,ip_9_29,p1270,p1271);
FA fa634(ip_10_28,ip_11_27,ip_12_26,p1272,p1273);
FA fa635(ip_13_25,ip_14_24,ip_15_23,p1274,p1275);
FA fa636(ip_16_22,ip_17_21,ip_18_20,p1276,p1277);
HA ha2(ip_19_19,ip_20_18,p1278,p1279);
FA fa637(ip_21_17,ip_22_16,ip_23_15,p1280,p1281);
FA fa638(ip_24_14,ip_25_13,ip_26_12,p1282,p1283);
FA fa639(ip_27_11,ip_28_10,ip_29_9,p1284,p1285);
FA fa640(ip_30_8,ip_31_7,p1279,p1286,p1287);
FA fa641(p1271,p1273,p1275,p1288,p1289);
FA fa642(p1277,p1281,p1283,p1290,p1291);
FA fa643(p1285,p1287,p1218,p1292,p1293);
FA fa644(p1220,p1222,p1224,p1294,p1295);
FA fa645(p1226,p1228,p1230,p1296,p1297);
FA fa646(p1232,p1234,p1289,p1298,p1299);
FA fa647(p1291,p1293,p1236,p1300,p1301);
FA fa648(p1238,p1295,p1297,p1302,p1303);
FA fa649(p1240,p1242,p1244,p1304,p1305);
HA ha3(p1246,p1299,p1306,p1307);
FA fa650(p1301,p1303,p1307,p1308,p1309);
FA fa651(p1248,p1250,p1252,p1310,p1311);
FA fa652(p1305,p1254,p1309,p1312,p1313);
FA fa653(p1256,p1311,p1258,p1314,p1315);
FA fa654(p1313,p1260,p1315,p1316,p1317);
FA fa655(p1262,p1317,p1264,p1318,p1319);
FA fa656(p1319,p1266,p1268,p1320,p1321);
FA fa657(ip_8_31,ip_9_30,ip_10_29,p1322,p1323);
FA fa658(ip_11_28,ip_12_27,ip_13_26,p1324,p1325);
FA fa659(ip_14_25,ip_15_24,ip_16_23,p1326,p1327);
FA fa660(ip_17_22,ip_18_21,ip_19_20,p1328,p1329);
FA fa661(ip_20_19,ip_21_18,ip_22_17,p1330,p1331);
FA fa662(ip_23_16,ip_24_15,ip_25_14,p1332,p1333);
FA fa663(ip_26_13,ip_27_12,ip_28_11,p1334,p1335);
FA fa664(ip_29_10,ip_30_9,ip_31_8,p1336,p1337);
FA fa665(p1278,p1323,p1325,p1338,p1339);
FA fa666(p1327,p1329,p1331,p1340,p1341);
FA fa667(p1333,p1335,p1337,p1342,p1343);
FA fa668(p1270,p1272,p1274,p1344,p1345);
FA fa669(p1276,p1280,p1282,p1346,p1347);
FA fa670(p1284,p1286,p1339,p1348,p1349);
FA fa671(p1341,p1343,p1288,p1350,p1351);
FA fa672(p1290,p1292,p1345,p1352,p1353);
FA fa673(p1347,p1349,p1294,p1354,p1355);
FA fa674(p1296,p1351,p1298,p1356,p1357);
FA fa675(p1300,p1306,p1353,p1358,p1359);
FA fa676(p1355,p1302,p1357,p1360,p1361);
FA fa677(p1304,p1359,p1308,p1362,p1363);
FA fa678(p1361,p1310,p1363,p1364,p1365);
FA fa679(p1312,p1314,p1365,p1366,p1367);
FA fa680(p1316,p1367,p1318,p1368,p1369);
FA fa681(ip_9_31,ip_10_30,ip_11_29,p1370,p1371);
FA fa682(ip_12_28,ip_13_27,ip_14_26,p1372,p1373);
FA fa683(ip_15_25,ip_16_24,ip_17_23,p1374,p1375);
FA fa684(ip_18_22,ip_19_21,ip_20_20,p1376,p1377);
FA fa685(ip_21_19,ip_22_18,ip_23_17,p1378,p1379);
FA fa686(ip_24_16,ip_25_15,ip_26_14,p1380,p1381);
FA fa687(ip_27_13,ip_28_12,ip_29_11,p1382,p1383);
FA fa688(ip_30_10,ip_31_9,p1371,p1384,p1385);
FA fa689(p1373,p1375,p1377,p1386,p1387);
FA fa690(p1379,p1381,p1383,p1388,p1389);
FA fa691(p1322,p1324,p1326,p1390,p1391);
FA fa692(p1328,p1330,p1332,p1392,p1393);
HA ha4(p1334,p1336,p1394,p1395);
FA fa693(p1385,p1387,p1389,p1396,p1397);
FA fa694(p1395,p1338,p1340,p1398,p1399);
FA fa695(p1342,p1391,p1393,p1400,p1401);
FA fa696(p1344,p1346,p1348,p1402,p1403);
FA fa697(p1397,p1350,p1399,p1404,p1405);
FA fa698(p1401,p1352,p1354,p1406,p1407);
FA fa699(p1403,p1356,p1405,p1408,p1409);
FA fa700(p1358,p1407,p1360,p1410,p1411);
FA fa701(p1409,p1362,p1411,p1412,p1413);
FA fa702(p1364,p1413,p1366,p1414,p1415);
FA fa703(ip_10_31,ip_11_30,ip_12_29,p1416,p1417);
HA ha5(ip_13_28,ip_14_27,p1418,p1419);
FA fa704(ip_15_26,ip_16_25,ip_17_24,p1420,p1421);
FA fa705(ip_18_23,ip_19_22,ip_20_21,p1422,p1423);
FA fa706(ip_21_20,ip_22_19,ip_23_18,p1424,p1425);
FA fa707(ip_24_17,ip_25_16,ip_26_15,p1426,p1427);
FA fa708(ip_27_14,ip_28_13,ip_29_12,p1428,p1429);
FA fa709(ip_30_11,ip_31_10,p1419,p1430,p1431);
FA fa710(p1417,p1421,p1423,p1432,p1433);
HA ha6(p1425,p1427,p1434,p1435);
FA fa711(p1429,p1431,p1370,p1436,p1437);
HA ha7(p1372,p1374,p1438,p1439);
FA fa712(p1376,p1378,p1380,p1440,p1441);
FA fa713(p1382,p1435,p1384,p1442,p1443);
HA ha8(p1394,p1433,p1444,p1445);
FA fa714(p1437,p1439,p1386,p1446,p1447);
FA fa715(p1388,p1441,p1443,p1448,p1449);
FA fa716(p1445,p1390,p1392,p1450,p1451);
FA fa717(p1447,p1396,p1449,p1452,p1453);
FA fa718(p1398,p1400,p1451,p1454,p1455);
FA fa719(p1402,p1453,p1404,p1456,p1457);
FA fa720(p1455,p1406,p1457,p1458,p1459);
FA fa721(p1408,p1410,p1459,p1460,p1461);
FA fa722(p1412,p1461,p1414,p1462,p1463);
FA fa723(ip_11_31,ip_12_30,ip_13_29,p1464,p1465);
FA fa724(ip_14_28,ip_15_27,ip_16_26,p1466,p1467);
FA fa725(ip_17_25,ip_18_24,ip_19_23,p1468,p1469);
FA fa726(ip_20_22,ip_21_21,ip_22_20,p1470,p1471);
FA fa727(ip_23_19,ip_24_18,ip_25_17,p1472,p1473);
FA fa728(ip_26_16,ip_27_15,ip_28_14,p1474,p1475);
FA fa729(ip_29_13,ip_30_12,ip_31_11,p1476,p1477);
FA fa730(p1418,p1465,p1467,p1478,p1479);
HA ha9(p1469,p1471,p1480,p1481);
HA ha10(p1473,p1475,p1482,p1483);
FA fa731(p1477,p1416,p1420,p1484,p1485);
FA fa732(p1422,p1424,p1426,p1486,p1487);
FA fa733(p1428,p1430,p1434,p1488,p1489);
FA fa734(p1481,p1483,p1438,p1490,p1491);
FA fa735(p1479,p1432,p1436,p1492,p1493);
FA fa736(p1444,p1485,p1487,p1494,p1495);
FA fa737(p1489,p1491,p1440,p1496,p1497);
FA fa738(p1442,p1446,p1493,p1498,p1499);
HA ha11(p1495,p1497,p1500,p1501);
FA fa739(p1448,p1501,p1450,p1502,p1503);
FA fa740(p1499,p1452,p1503,p1504,p1505);
HA ha12(p1454,p1456,p1506,p1507);
FA fa741(p1505,p1507,p1458,p1508,p1509);
FA fa742(p1509,p1460,p1462,p1510,p1511);
FA fa743(ip_12_31,ip_13_30,ip_14_29,p1512,p1513);
HA ha13(ip_15_28,ip_16_27,p1514,p1515);
FA fa744(ip_17_26,ip_18_25,ip_19_24,p1516,p1517);
FA fa745(ip_20_23,ip_21_22,ip_22_21,p1518,p1519);
FA fa746(ip_23_20,ip_24_19,ip_25_18,p1520,p1521);
HA ha14(ip_26_17,ip_27_16,p1522,p1523);
FA fa747(ip_28_15,ip_29_14,ip_30_13,p1524,p1525);
FA fa748(ip_31_12,p1515,p1523,p1526,p1527);
FA fa749(p1513,p1517,p1519,p1528,p1529);
FA fa750(p1521,p1525,p1464,p1530,p1531);
FA fa751(p1466,p1468,p1470,p1532,p1533);
FA fa752(p1472,p1474,p1476,p1534,p1535);
FA fa753(p1480,p1482,p1527,p1536,p1537);
FA fa754(p1529,p1531,p1478,p1538,p1539);
FA fa755(p1533,p1535,p1537,p1540,p1541);
FA fa756(p1484,p1486,p1488,p1542,p1543);
FA fa757(p1490,p1539,p1541,p1544,p1545);
FA fa758(p1492,p1494,p1496,p1546,p1547);
FA fa759(p1500,p1543,p1545,p1548,p1549);
FA fa760(p1498,p1547,p1549,p1550,p1551);
HA ha15(p1502,p1551,p1552,p1553);
FA fa761(p1504,p1506,p1553,p1554,p1555);
FA fa762(p1555,p1508,p1510,p1556,p1557);
FA fa763(ip_13_31,ip_14_30,ip_15_29,p1558,p1559);
FA fa764(ip_16_28,ip_17_27,ip_18_26,p1560,p1561);
FA fa765(ip_19_25,ip_20_24,ip_21_23,p1562,p1563);
FA fa766(ip_22_22,ip_23_21,ip_24_20,p1564,p1565);
FA fa767(ip_25_19,ip_26_18,ip_27_17,p1566,p1567);
FA fa768(ip_28_16,ip_29_15,ip_30_14,p1568,p1569);
FA fa769(ip_31_13,p1514,p1522,p1570,p1571);
FA fa770(p1559,p1561,p1563,p1572,p1573);
FA fa771(p1565,p1567,p1569,p1574,p1575);
FA fa772(p1512,p1516,p1518,p1576,p1577);
FA fa773(p1520,p1524,p1571,p1578,p1579);
FA fa774(p1526,p1573,p1575,p1580,p1581);
FA fa775(p1528,p1530,p1577,p1582,p1583);
FA fa776(p1579,p1532,p1534,p1584,p1585);
FA fa777(p1536,p1581,p1538,p1586,p1587);
HA ha16(p1583,p1540,p1588,p1589);
FA fa778(p1585,p1587,p1542,p1590,p1591);
HA ha17(p1544,p1589,p1592,p1593);
FA fa779(p1591,p1593,p1546,p1594,p1595);
FA fa780(p1548,p1595,p1550,p1596,p1597);
FA fa781(p1552,p1597,p1554,p1598,p1599);
FA fa782(ip_14_31,ip_15_30,ip_16_29,p1600,p1601);
FA fa783(ip_17_28,ip_18_27,ip_19_26,p1602,p1603);
HA ha18(ip_20_25,ip_21_24,p1604,p1605);
HA ha19(ip_22_23,ip_23_22,p1606,p1607);
FA fa784(ip_24_21,ip_25_20,ip_26_19,p1608,p1609);
FA fa785(ip_27_18,ip_28_17,ip_29_16,p1610,p1611);
FA fa786(ip_30_15,ip_31_14,p1605,p1612,p1613);
FA fa787(p1607,p1601,p1603,p1614,p1615);
FA fa788(p1609,p1611,p1613,p1616,p1617);
HA ha20(p1558,p1560,p1618,p1619);
FA fa789(p1562,p1564,p1566,p1620,p1621);
HA ha21(p1568,p1570,p1622,p1623);
FA fa790(p1615,p1617,p1619,p1624,p1625);
FA fa791(p1572,p1574,p1621,p1626,p1627);
FA fa792(p1623,p1576,p1578,p1628,p1629);
HA ha22(p1625,p1580,p1630,p1631);
FA fa793(p1627,p1582,p1629,p1632,p1633);
FA fa794(p1631,p1584,p1586,p1634,p1635);
FA fa795(p1588,p1592,p1633,p1636,p1637);
FA fa796(p1590,p1635,p1637,p1638,p1639);
FA fa797(p1594,p1639,p1596,p1640,p1641);
FA fa798(ip_15_31,ip_16_30,ip_17_29,p1642,p1643);
FA fa799(ip_18_28,ip_19_27,ip_20_26,p1644,p1645);
HA ha23(ip_21_25,ip_22_24,p1646,p1647);
FA fa800(ip_23_23,ip_24_22,ip_25_21,p1648,p1649);
HA ha24(ip_26_20,ip_27_19,p1650,p1651);
FA fa801(ip_28_18,ip_29_17,ip_30_16,p1652,p1653);
FA fa802(ip_31_15,p1604,p1606,p1654,p1655);
FA fa803(p1647,p1651,p1643,p1656,p1657);
HA ha25(p1645,p1649,p1658,p1659);
FA fa804(p1653,p1600,p1602,p1660,p1661);
FA fa805(p1608,p1610,p1612,p1662,p1663);
FA fa806(p1655,p1657,p1659,p1664,p1665);
FA fa807(p1618,p1614,p1616,p1666,p1667);
FA fa808(p1622,p1661,p1663,p1668,p1669);
FA fa809(p1665,p1620,p1624,p1670,p1671);
FA fa810(p1667,p1669,p1626,p1672,p1673);
HA ha26(p1630,p1671,p1674,p1675);
FA fa811(p1628,p1673,p1675,p1676,p1677);
HA ha27(p1632,p1677,p1678,p1679);
HA ha28(p1634,p1679,p1680,p1681);
FA fa812(p1636,p1681,p1638,p1682,p1683);
FA fa813(ip_16_31,ip_17_30,ip_18_29,p1684,p1685);
FA fa814(ip_19_28,ip_20_27,ip_21_26,p1686,p1687);
HA ha29(ip_22_25,ip_23_24,p1688,p1689);
FA fa815(ip_24_23,ip_25_22,ip_26_21,p1690,p1691);
FA fa816(ip_27_20,ip_28_19,ip_29_18,p1692,p1693);
HA ha30(ip_30_17,ip_31_16,p1694,p1695);
HA ha31(p1646,p1650,p1696,p1697);
HA ha32(p1689,p1695,p1698,p1699);
HA ha33(p1685,p1687,p1700,p1701);
FA fa817(p1691,p1693,p1697,p1702,p1703);
HA ha34(p1699,p1642,p1704,p1705);
FA fa818(p1644,p1648,p1652,p1706,p1707);
HA ha35(p1658,p1701,p1708,p1709);
FA fa819(p1654,p1656,p1703,p1710,p1711);
FA fa820(p1705,p1709,p1707,p1712,p1713);
FA fa821(p1660,p1662,p1664,p1714,p1715);
FA fa822(p1711,p1713,p1666,p1716,p1717);
HA ha36(p1668,p1715,p1718,p1719);
FA fa823(p1670,p1674,p1717,p1720,p1721);
FA fa824(p1719,p1672,p1721,p1722,p1723);
HA ha37(p1676,p1678,p1724,p1725);
HA ha38(p1723,p1680,p1726,p1727);
FA fa825(p1725,p1727,p1682,p1728,p1729);
HA ha39(ip_17_31,ip_18_30,p1730,p1731);
FA fa826(ip_19_29,ip_20_28,ip_21_27,p1732,p1733);
FA fa827(ip_22_26,ip_23_25,ip_24_24,p1734,p1735);
FA fa828(ip_25_23,ip_26_22,ip_27_21,p1736,p1737);
HA ha40(ip_28_20,ip_29_19,p1738,p1739);
FA fa829(ip_30_18,ip_31_17,p1688,p1740,p1741);
FA fa830(p1694,p1731,p1739,p1742,p1743);
FA fa831(p1696,p1698,p1733,p1744,p1745);
FA fa832(p1735,p1737,p1741,p1746,p1747);
HA ha41(p1684,p1686,p1748,p1749);
FA fa833(p1690,p1692,p1700,p1750,p1751);
FA fa834(p1743,p1704,p1708,p1752,p1753);
FA fa835(p1745,p1747,p1749,p1754,p1755);
HA ha42(p1702,p1751,p1756,p1757);
HA ha43(p1706,p1753,p1758,p1759);
FA fa836(p1755,p1757,p1710,p1760,p1761);
FA fa837(p1712,p1759,p1761,p1762,p1763);
HA ha44(p1714,p1718,p1764,p1765);
HA ha45(p1763,p1716,p1766,p1767);
HA ha46(p1765,p1767,p1768,p1769);
FA fa838(p1720,p1769,p1722,p1770,p1771);
FA fa839(p1724,p1726,p1771,p1772,p1773);
HA ha47(ip_18_31,ip_19_30,p1774,p1775);
FA fa840(ip_20_29,ip_21_28,ip_22_27,p1776,p1777);
HA ha48(ip_23_26,ip_24_25,p1778,p1779);
HA ha49(ip_25_24,ip_26_23,p1780,p1781);
HA ha50(ip_27_22,ip_28_21,p1782,p1783);
FA fa841(ip_29_20,ip_30_19,ip_31_18,p1784,p1785);
HA ha51(p1730,p1738,p1786,p1787);
FA fa842(p1775,p1779,p1781,p1788,p1789);
HA ha52(p1783,p1777,p1790,p1791);
HA ha53(p1785,p1787,p1792,p1793);
HA ha54(p1732,p1734,p1794,p1795);
FA fa843(p1736,p1740,p1789,p1796,p1797);
HA ha55(p1791,p1793,p1798,p1799);
FA fa844(p1742,p1748,p1795,p1800,p1801);
HA ha56(p1799,p1744,p1802,p1803);
HA ha57(p1746,p1797,p1804,p1805);
FA fa845(p1750,p1756,p1801,p1806,p1807);
HA ha58(p1803,p1805,p1808,p1809);
HA ha59(p1752,p1754,p1810,p1811);
HA ha60(p1758,p1809,p1812,p1813);
HA ha61(p1807,p1811,p1814,p1815);
HA ha62(p1813,p1760,p1816,p1817);
HA ha63(p1815,p1762,p1818,p1819);
FA fa846(p1764,p1817,p1766,p1820,p1821);
HA ha64(p1819,p1768,p1822,p1823);
FA fa847(p1821,p1823,p1770,p1824,p1825);
HA ha65(ip_19_31,ip_20_30,p1826,p1827);
HA ha66(ip_21_29,ip_22_28,p1828,p1829);
FA fa848(ip_23_27,ip_24_26,ip_25_25,p1830,p1831);
HA ha67(ip_26_24,ip_27_23,p1832,p1833);
HA ha68(ip_28_22,ip_29_21,p1834,p1835);
HA ha69(ip_30_20,ip_31_19,p1836,p1837);
FA fa849(p1774,p1778,p1780,p1838,p1839);
HA ha70(p1782,p1827,p1840,p1841);
HA ha71(p1829,p1833,p1842,p1843);
HA ha72(p1835,p1837,p1844,p1845);
FA fa850(p1786,p1831,p1841,p1846,p1847);
FA fa851(p1843,p1845,p1776,p1848,p1849);
HA ha73(p1784,p1790,p1850,p1851);
HA ha74(p1792,p1839,p1852,p1853);
HA ha75(p1788,p1794,p1854,p1855);
FA fa852(p1798,p1847,p1849,p1856,p1857);
HA ha76(p1851,p1853,p1858,p1859);
HA ha77(p1855,p1859,p1860,p1861);
FA fa853(p1796,p1802,p1804,p1862,p1863);
HA ha78(p1857,p1861,p1864,p1865);
HA ha79(p1800,p1808,p1866,p1867);
HA ha80(p1865,p1810,p1868,p1869);
FA fa854(p1812,p1863,p1867,p1870,p1871);
HA ha81(p1806,p1814,p1872,p1873);
HA ha82(p1869,p1816,p1874,p1875);
HA ha83(p1871,p1873,p1876,p1877);
FA fa855(p1818,p1875,p1877,p1878,p1879);
FA fa856(p1820,p1822,p1879,p1880,p1881);
FA fa857(ip_20_31,ip_21_30,ip_22_29,p1882,p1883);
FA fa858(ip_23_28,ip_24_27,ip_25_26,p1884,p1885);
HA ha84(ip_26_25,ip_27_24,p1886,p1887);
HA ha85(ip_28_23,ip_29_22,p1888,p1889);
HA ha86(ip_30_21,ip_31_20,p1890,p1891);
FA fa859(p1826,p1828,p1832,p1892,p1893);
HA ha87(p1834,p1836,p1894,p1895);
HA ha88(p1887,p1889,p1896,p1897);
FA fa860(p1891,p1840,p1842,p1898,p1899);
HA ha89(p1844,p1883,p1900,p1901);
HA ha90(p1885,p1895,p1902,p1903);
HA ha91(p1897,p1830,p1904,p1905);
HA ha92(p1893,p1901,p1906,p1907);
HA ha93(p1903,p1838,p1908,p1909);
HA ha94(p1850,p1852,p1910,p1911);
HA ha95(p1899,p1905,p1912,p1913);
HA ha96(p1907,p1846,p1914,p1915);
FA fa861(p1848,p1854,p1858,p1916,p1917);
HA ha97(p1909,p1911,p1918,p1919);
FA fa862(p1913,p1860,p1915,p1920,p1921);
HA ha98(p1919,p1856,p1922,p1923);
HA ha99(p1864,p1917,p1924,p1925);
HA ha100(p1866,p1921,p1926,p1927);
HA ha101(p1923,p1925,p1928,p1929);
HA ha102(p1862,p1868,p1930,p1931);
HA ha103(p1927,p1929,p1932,p1933);
HA ha104(p1872,p1931,p1934,p1935);
HA ha105(p1933,p1870,p1936,p1937);
HA ha106(p1874,p1876,p1938,p1939);
FA fa863(p1935,p1937,p1939,p1940,p1941);
HA ha107(p1878,p1941,p1942,p1943);
FA fa864(ip_21_31,ip_22_30,ip_23_29,p1944,p1945);
FA fa865(ip_24_28,ip_25_27,ip_26_26,p1946,p1947);
HA ha108(ip_27_25,ip_28_24,p1948,p1949);
HA ha109(ip_29_23,ip_30_22,p1950,p1951);
HA ha110(ip_31_21,p1886,p1952,p1953);
FA fa866(p1888,p1890,p1949,p1954,p1955);
FA fa867(p1951,p1894,p1896,p1956,p1957);
HA ha111(p1945,p1947,p1958,p1959);
HA ha112(p1953,p1882,p1960,p1961);
HA ha113(p1884,p1900,p1962,p1963);
HA ha114(p1902,p1955,p1964,p1965);
FA fa868(p1959,p1892,p1904,p1966,p1967);
HA ha115(p1906,p1957,p1968,p1969);
FA fa869(p1961,p1963,p1965,p1970,p1971);
FA fa870(p1898,p1908,p1910,p1972,p1973);
HA ha116(p1912,p1969,p1974,p1975);
HA ha117(p1914,p1918,p1976,p1977);
HA ha118(p1967,p1971,p1978,p1979);
HA ha119(p1975,p1973,p1980,p1981);
HA ha120(p1977,p1979,p1982,p1983);
HA ha121(p1916,p1922,p1984,p1985);
FA fa871(p1924,p1981,p1983,p1986,p1987);
HA ha122(p1920,p1926,p1988,p1989);
HA ha123(p1928,p1985,p1990,p1991);
FA fa872(p1930,p1932,p1987,p1992,p1993);
HA ha124(p1989,p1991,p1994,p1995);
HA ha125(p1934,p1995,p1996,p1997);
HA ha126(p1936,p1938,p1998,p1999);
HA ha127(p1993,p1997,p2000,p2001);
HA ha128(p1999,p2001,p2002,p2003);
HA ha129(p2003,p1940,p2004,p2005);
HA ha130(ip_22_31,ip_23_30,p2006,p2007);
HA ha131(ip_24_29,ip_25_28,p2008,p2009);
HA ha132(ip_26_27,ip_27_26,p2010,p2011);
HA ha133(ip_28_25,ip_29_24,p2012,p2013);
HA ha134(ip_30_23,ip_31_22,p2014,p2015);
FA fa873(p1948,p1950,p2007,p2016,p2017);
HA ha135(p2009,p2011,p2018,p2019);
HA ha136(p2013,p2015,p2020,p2021);
HA ha137(p1952,p2019,p2022,p2023);
HA ha138(p2021,p1944,p2024,p2025);
HA ha139(p1946,p1958,p2026,p2027);
HA ha140(p2017,p2023,p2028,p2029);
HA ha141(p1954,p1960,p2030,p2031);
HA ha142(p1962,p1964,p2032,p2033);
HA ha143(p2025,p2027,p2034,p2035);
HA ha144(p2029,p1956,p2036,p2037);
HA ha145(p1968,p2031,p2038,p2039);
HA ha146(p2033,p2035,p2040,p2041);
HA ha147(p1974,p2037,p2042,p2043);
HA ha148(p2039,p2041,p2044,p2045);
HA ha149(p1966,p1970,p2046,p2047);
HA ha150(p1976,p1978,p2048,p2049);
HA ha151(p2043,p2045,p2050,p2051);
HA ha152(p1972,p1980,p2052,p2053);
HA ha153(p1982,p2047,p2054,p2055);
FA fa874(p2049,p2051,p1984,p2056,p2057);
FA fa875(p2053,p2055,p1988,p2058,p2059);
HA ha154(p1990,p2057,p2060,p2061);
HA ha155(p1986,p1994,p2062,p2063);
HA ha156(p2059,p2061,p2064,p2065);
HA ha157(p1996,p2063,p2066,p2067);
HA ha158(p2065,p1992,p2068,p2069);
HA ha159(p1998,p2000,p2070,p2071);
HA ha160(p2067,p2002,p2072,p2073);
HA ha161(p2069,p2071,p2074,p2075);
HA ha162(p2073,p2075,p2076,p2077);
HA ha163(ip_23_31,ip_24_30,p2078,p2079);
HA ha164(ip_25_29,ip_26_28,p2080,p2081);
HA ha165(ip_27_27,ip_28_26,p2082,p2083);
HA ha166(ip_29_25,ip_30_24,p2084,p2085);
HA ha167(ip_31_23,p2006,p2086,p2087);
FA fa876(p2008,p2010,p2012,p2088,p2089);
HA ha168(p2014,p2079,p2090,p2091);
HA ha169(p2081,p2083,p2092,p2093);
FA fa877(p2085,p2018,p2020,p2094,p2095);
HA ha170(p2087,p2091,p2096,p2097);
HA ha171(p2093,p2022,p2098,p2099);
HA ha172(p2089,p2097,p2100,p2101);
HA ha173(p2016,p2024,p2102,p2103);
HA ha174(p2026,p2028,p2104,p2105);
HA ha175(p2095,p2099,p2106,p2107);
HA ha176(p2101,p2030,p2108,p2109);
FA fa878(p2032,p2034,p2103,p2110,p2111);
HA ha177(p2105,p2107,p2112,p2113);
HA ha178(p2036,p2038,p2114,p2115);
HA ha179(p2040,p2109,p2116,p2117);
HA ha180(p2113,p2042,p2118,p2119);
HA ha181(p2044,p2111,p2120,p2121);
HA ha182(p2115,p2117,p2122,p2123);
HA ha183(p2046,p2048,p2124,p2125);
HA ha184(p2050,p2119,p2126,p2127);
HA ha185(p2121,p2123,p2128,p2129);
FA fa879(p2052,p2054,p2125,p2130,p2131);
HA ha186(p2127,p2129,p2132,p2133);
HA ha187(p2133,p2056,p2134,p2135);
HA ha188(p2060,p2131,p2136,p2137);
HA ha189(p2058,p2062,p2138,p2139);
HA ha190(p2064,p2135,p2140,p2141);
HA ha191(p2137,p2066,p2142,p2143);
HA ha192(p2139,p2141,p2144,p2145);
FA fa880(p2068,p2070,p2143,p2146,p2147);
HA ha193(p2145,p2072,p2148,p2149);
HA ha194(p2074,p2076,p2150,p2151);
HA ha195(p2147,p2149,p2152,p2153);
HA ha196(ip_24_31,ip_25_30,p2154,p2155);
HA ha197(ip_26_29,ip_27_28,p2156,p2157);
HA ha198(ip_28_27,ip_29_26,p2158,p2159);
HA ha199(ip_30_25,ip_31_24,p2160,p2161);
HA ha200(p2078,p2080,p2162,p2163);
HA ha201(p2082,p2084,p2164,p2165);
HA ha202(p2155,p2157,p2166,p2167);
HA ha203(p2159,p2161,p2168,p2169);
HA ha204(p2086,p2090,p2170,p2171);
HA ha205(p2092,p2163,p2172,p2173);
HA ha206(p2165,p2167,p2174,p2175);
HA ha207(p2169,p2096,p2176,p2177);
HA ha208(p2171,p2173,p2178,p2179);
HA ha209(p2175,p2088,p2180,p2181);
HA ha210(p2098,p2100,p2182,p2183);
HA ha211(p2177,p2179,p2184,p2185);
HA ha212(p2094,p2102,p2186,p2187);
HA ha213(p2104,p2106,p2188,p2189);
HA ha214(p2181,p2183,p2190,p2191);
HA ha215(p2185,p2108,p2192,p2193);
HA ha216(p2112,p2187,p2194,p2195);
HA ha217(p2189,p2191,p2196,p2197);
HA ha218(p2114,p2116,p2198,p2199);
HA ha219(p2193,p2195,p2200,p2201);
HA ha220(p2197,p2110,p2202,p2203);
HA ha221(p2118,p2120,p2204,p2205);
HA ha222(p2122,p2199,p2206,p2207);
HA ha223(p2201,p2124,p2208,p2209);
HA ha224(p2126,p2128,p2210,p2211);
HA ha225(p2203,p2205,p2212,p2213);
HA ha226(p2207,p2132,p2214,p2215);
HA ha227(p2209,p2211,p2216,p2217);
HA ha228(p2213,p2215,p2218,p2219);
HA ha229(p2217,p2130,p2220,p2221);
HA ha230(p2134,p2136,p2222,p2223);
HA ha231(p2219,p2138,p2224,p2225);
HA ha232(p2140,p2221,p2226,p2227);
HA ha233(p2223,p2142,p2228,p2229);
HA ha234(p2144,p2225,p2230,p2231);
HA ha235(p2227,p2229,p2232,p2233);
HA ha236(p2231,p2148,p2234,p2235);
HA ha237(p2233,p2146,p2236,p2237);
HA ha238(p2150,p2152,p2238,p2239);
HA ha239(p2235,p2237,p2240,p2241);
HA ha240(ip_25_31,ip_26_30,p2242,p2243);
HA ha241(ip_27_29,ip_28_28,p2244,p2245);
HA ha242(ip_29_27,ip_30_26,p2246,p2247);
HA ha243(ip_31_25,p2154,p2248,p2249);
HA ha244(p2156,p2158,p2250,p2251);
HA ha245(p2160,p2243,p2252,p2253);
HA ha246(p2245,p2247,p2254,p2255);
HA ha247(p2162,p2164,p2256,p2257);
HA ha248(p2166,p2168,p2258,p2259);
HA ha249(p2249,p2251,p2260,p2261);
HA ha250(p2253,p2255,p2262,p2263);
HA ha251(p2170,p2172,p2264,p2265);
HA ha252(p2174,p2257,p2266,p2267);
HA ha253(p2259,p2261,p2268,p2269);
HA ha254(p2263,p2176,p2270,p2271);
HA ha255(p2178,p2265,p2272,p2273);
HA ha256(p2267,p2269,p2274,p2275);
FA fa881(p2180,p2182,p2184,p2276,p2277);
HA ha257(p2271,p2273,p2278,p2279);
HA ha258(p2275,p2186,p2280,p2281);
HA ha259(p2188,p2190,p2282,p2283);
HA ha260(p2279,p2192,p2284,p2285);
HA ha261(p2194,p2196,p2286,p2287);
HA ha262(p2277,p2281,p2288,p2289);
HA ha263(p2283,p2198,p2290,p2291);
FA fa882(p2200,p2285,p2287,p2292,p2293);
HA ha264(p2289,p2202,p2294,p2295);
HA ha265(p2204,p2206,p2296,p2297);
FA fa883(p2291,p2208,p2210,p2298,p2299);
HA ha266(p2212,p2293,p2300,p2301);
HA ha267(p2295,p2297,p2302,p2303);
HA ha268(p2214,p2216,p2304,p2305);
HA ha269(p2301,p2303,p2306,p2307);
HA ha270(p2218,p2299,p2308,p2309);
FA fa884(p2305,p2307,p2220,p2310,p2311);
HA ha271(p2222,p2309,p2312,p2313);
HA ha272(p2224,p2226,p2314,p2315);
HA ha273(p2311,p2313,p2316,p2317);
HA ha274(p2228,p2230,p2318,p2319);
HA ha275(p2315,p2317,p2320,p2321);
HA ha276(p2232,p2319,p2322,p2323);
HA ha277(p2321,p2234,p2324,p2325);
FA fa885(p2323,p2236,p2238,p2326,p2327);
HA ha278(p2325,p2240,p2328,p2329);
HA ha279(ip_26_31,ip_27_30,p2330,p2331);
HA ha280(ip_28_29,ip_29_28,p2332,p2333);
HA ha281(ip_30_27,ip_31_26,p2334,p2335);
HA ha282(p2242,p2244,p2336,p2337);
HA ha283(p2246,p2331,p2338,p2339);
FA fa886(p2333,p2335,p2248,p2340,p2341);
HA ha284(p2250,p2252,p2342,p2343);
HA ha285(p2254,p2337,p2344,p2345);
HA ha286(p2339,p2256,p2346,p2347);
HA ha287(p2258,p2260,p2348,p2349);
HA ha288(p2262,p2341,p2350,p2351);
HA ha289(p2343,p2345,p2352,p2353);
HA ha290(p2264,p2266,p2354,p2355);
HA ha291(p2268,p2347,p2356,p2357);
HA ha292(p2349,p2351,p2358,p2359);
HA ha293(p2353,p2270,p2360,p2361);
HA ha294(p2272,p2274,p2362,p2363);
HA ha295(p2355,p2357,p2364,p2365);
HA ha296(p2359,p2278,p2366,p2367);
HA ha297(p2361,p2363,p2368,p2369);
HA ha298(p2365,p2280,p2370,p2371);
HA ha299(p2282,p2367,p2372,p2373);
HA ha300(p2369,p2276,p2374,p2375);
HA ha301(p2284,p2286,p2376,p2377);
HA ha302(p2288,p2371,p2378,p2379);
HA ha303(p2373,p2290,p2380,p2381);
HA ha304(p2375,p2377,p2382,p2383);
HA ha305(p2379,p2294,p2384,p2385);
HA ha306(p2296,p2381,p2386,p2387);
HA ha307(p2383,p2292,p2388,p2389);
HA ha308(p2300,p2302,p2390,p2391);
HA ha309(p2385,p2387,p2392,p2393);
HA ha310(p2304,p2306,p2394,p2395);
HA ha311(p2389,p2391,p2396,p2397);
HA ha312(p2393,p2298,p2398,p2399);
HA ha313(p2308,p2395,p2400,p2401);
HA ha314(p2397,p2312,p2402,p2403);
HA ha315(p2399,p2401,p2404,p2405);
HA ha316(p2310,p2314,p2406,p2407);
HA ha317(p2316,p2403,p2408,p2409);
HA ha318(p2405,p2318,p2410,p2411);
HA ha319(p2320,p2407,p2412,p2413);
HA ha320(p2409,p2322,p2414,p2415);
HA ha321(p2411,p2413,p2416,p2417);
HA ha322(p2324,p2415,p2418,p2419);
HA ha323(p2417,p2419,p2420,p2421);
HA ha324(p2328,p2421,p2422,p2423);
HA ha325(ip_27_31,ip_28_30,p2424,p2425);
HA ha326(ip_29_29,ip_30_28,p2426,p2427);
HA ha327(ip_31_27,p2330,p2428,p2429);
HA ha328(p2332,p2334,p2430,p2431);
HA ha329(p2425,p2427,p2432,p2433);
HA ha330(p2336,p2338,p2434,p2435);
HA ha331(p2429,p2431,p2436,p2437);
HA ha332(p2433,p2342,p2438,p2439);
HA ha333(p2344,p2435,p2440,p2441);
HA ha334(p2437,p2340,p2442,p2443);
HA ha335(p2346,p2348,p2444,p2445);
HA ha336(p2350,p2352,p2446,p2447);
HA ha337(p2439,p2441,p2448,p2449);
HA ha338(p2354,p2356,p2450,p2451);
HA ha339(p2358,p2443,p2452,p2453);
HA ha340(p2445,p2447,p2454,p2455);
HA ha341(p2449,p2360,p2456,p2457);
HA ha342(p2362,p2364,p2458,p2459);
HA ha343(p2451,p2453,p2460,p2461);
HA ha344(p2455,p2366,p2462,p2463);
FA fa887(p2368,p2457,p2459,p2464,p2465);
HA ha345(p2461,p2370,p2466,p2467);
FA fa888(p2372,p2463,p2374,p2468,p2469);
FA fa889(p2376,p2378,p2465,p2470,p2471);
HA ha346(p2467,p2380,p2472,p2473);
HA ha347(p2382,p2469,p2474,p2475);
HA ha348(p2384,p2386,p2476,p2477);
HA ha349(p2471,p2473,p2478,p2479);
HA ha350(p2475,p2388,p2480,p2481);
HA ha351(p2390,p2392,p2482,p2483);
HA ha352(p2477,p2479,p2484,p2485);
HA ha353(p2394,p2396,p2486,p2487);
HA ha354(p2481,p2483,p2488,p2489);
HA ha355(p2485,p2398,p2490,p2491);
HA ha356(p2400,p2487,p2492,p2493);
HA ha357(p2489,p2402,p2494,p2495);
HA ha358(p2404,p2491,p2496,p2497);
HA ha359(p2493,p2406,p2498,p2499);
HA ha360(p2408,p2495,p2500,p2501);
HA ha361(p2497,p2410,p2502,p2503);
HA ha362(p2412,p2499,p2504,p2505);
HA ha363(p2501,p2414,p2506,p2507);
HA ha364(p2416,p2503,p2508,p2509);
HA ha365(p2505,p2418,p2510,p2511);
HA ha366(p2507,p2509,p2512,p2513);
HA ha367(p2420,p2511,p2514,p2515);
HA ha368(p2513,p2422,p2516,p2517);
HA ha369(ip_28_31,ip_29_30,p2518,p2519);
HA ha370(ip_30_29,ip_31_28,p2520,p2521);
HA ha371(p2424,p2426,p2522,p2523);
HA ha372(p2519,p2521,p2524,p2525);
HA ha373(p2428,p2430,p2526,p2527);
HA ha374(p2432,p2523,p2528,p2529);
HA ha375(p2525,p2434,p2530,p2531);
HA ha376(p2436,p2527,p2532,p2533);
HA ha377(p2529,p2438,p2534,p2535);
HA ha378(p2440,p2531,p2536,p2537);
HA ha379(p2533,p2442,p2538,p2539);
HA ha380(p2444,p2446,p2540,p2541);
HA ha381(p2448,p2535,p2542,p2543);
HA ha382(p2537,p2450,p2544,p2545);
HA ha383(p2452,p2454,p2546,p2547);
HA ha384(p2539,p2541,p2548,p2549);
HA ha385(p2543,p2456,p2550,p2551);
HA ha386(p2458,p2460,p2552,p2553);
HA ha387(p2545,p2547,p2554,p2555);
HA ha388(p2549,p2462,p2556,p2557);
HA ha389(p2551,p2553,p2558,p2559);
HA ha390(p2555,p2466,p2560,p2561);
HA ha391(p2557,p2559,p2562,p2563);
HA ha392(p2464,p2561,p2564,p2565);
HA ha393(p2563,p2468,p2566,p2567);
HA ha394(p2472,p2474,p2568,p2569);
HA ha395(p2565,p2470,p2570,p2571);
HA ha396(p2476,p2478,p2572,p2573);
HA ha397(p2567,p2569,p2574,p2575);
HA ha398(p2480,p2482,p2576,p2577);
HA ha399(p2484,p2571,p2578,p2579);
HA ha400(p2573,p2575,p2580,p2581);
HA ha401(p2486,p2488,p2582,p2583);
FA fa890(p2577,p2579,p2581,p2584,p2585);
HA ha402(p2490,p2492,p2586,p2587);
HA ha403(p2583,p2494,p2588,p2589);
HA ha404(p2496,p2585,p2590,p2591);
HA ha405(p2587,p2498,p2592,p2593);
HA ha406(p2500,p2589,p2594,p2595);
HA ha407(p2591,p2502,p2596,p2597);
HA ha408(p2504,p2593,p2598,p2599);
HA ha409(p2595,p2506,p2600,p2601);
HA ha410(p2508,p2597,p2602,p2603);
HA ha411(p2599,p2510,p2604,p2605);
HA ha412(p2512,p2601,p2606,p2607);
FA fa891(p2603,p2514,p2605,p2608,p2609);
HA ha413(p2607,p2516,p2610,p2611);
HA ha414(ip_29_31,ip_30_30,p2612,p2613);
HA ha415(ip_31_29,p2518,p2614,p2615);
HA ha416(p2520,p2613,p2616,p2617);
HA ha417(p2522,p2524,p2618,p2619);
HA ha418(p2615,p2617,p2620,p2621);
HA ha419(p2526,p2528,p2622,p2623);
HA ha420(p2619,p2621,p2624,p2625);
HA ha421(p2530,p2532,p2626,p2627);
HA ha422(p2623,p2625,p2628,p2629);
HA ha423(p2534,p2536,p2630,p2631);
HA ha424(p2627,p2629,p2632,p2633);
HA ha425(p2538,p2540,p2634,p2635);
HA ha426(p2542,p2631,p2636,p2637);
HA ha427(p2633,p2544,p2638,p2639);
HA ha428(p2546,p2548,p2640,p2641);
HA ha429(p2635,p2637,p2642,p2643);
HA ha430(p2550,p2552,p2644,p2645);
HA ha431(p2554,p2639,p2646,p2647);
HA ha432(p2641,p2643,p2648,p2649);
HA ha433(p2556,p2558,p2650,p2651);
HA ha434(p2645,p2647,p2652,p2653);
HA ha435(p2649,p2560,p2654,p2655);
HA ha436(p2562,p2651,p2656,p2657);
HA ha437(p2653,p2564,p2658,p2659);
HA ha438(p2655,p2657,p2660,p2661);
HA ha439(p2566,p2568,p2662,p2663);
HA ha440(p2659,p2661,p2664,p2665);
HA ha441(p2570,p2572,p2666,p2667);
HA ha442(p2574,p2663,p2668,p2669);
FA fa892(p2665,p2576,p2578,p2670,p2671);
HA ha443(p2580,p2667,p2672,p2673);
HA ha444(p2669,p2582,p2674,p2675);
HA ha445(p2673,p2586,p2676,p2677);
HA ha446(p2671,p2675,p2678,p2679);
HA ha447(p2584,p2588,p2680,p2681);
HA ha448(p2590,p2677,p2682,p2683);
HA ha449(p2679,p2592,p2684,p2685);
HA ha450(p2594,p2681,p2686,p2687);
HA ha451(p2683,p2596,p2688,p2689);
HA ha452(p2598,p2685,p2690,p2691);
HA ha453(p2687,p2600,p2692,p2693);
HA ha454(p2602,p2689,p2694,p2695);
HA ha455(p2691,p2604,p2696,p2697);
HA ha456(p2606,p2693,p2698,p2699);
HA ha457(p2695,p2697,p2700,p2701);
HA ha458(p2699,p2610,p2702,p2703);
HA ha459(p2701,p2608,p2704,p2705);
HA ha460(ip_30_31,ip_31_30,p2706,p2707);
HA ha461(p2612,p2707,p2708,p2709);
HA ha462(p2614,p2616,p2710,p2711);
HA ha463(p2709,p2618,p2712,p2713);
HA ha464(p2620,p2711,p2714,p2715);
HA ha465(p2622,p2624,p2716,p2717);
HA ha466(p2713,p2715,p2718,p2719);
FA fa893(p2626,p2628,p2717,p2720,p2721);
HA ha467(p2719,p2630,p2722,p2723);
HA ha468(p2632,p2634,p2724,p2725);
HA ha469(p2636,p2721,p2726,p2727);
HA ha470(p2723,p2638,p2728,p2729);
HA ha471(p2640,p2642,p2730,p2731);
HA ha472(p2725,p2727,p2732,p2733);
HA ha473(p2644,p2646,p2734,p2735);
HA ha474(p2648,p2729,p2736,p2737);
FA fa894(p2731,p2733,p2650,p2738,p2739);
HA ha475(p2652,p2735,p2740,p2741);
HA ha476(p2737,p2654,p2742,p2743);
HA ha477(p2656,p2739,p2744,p2745);
HA ha478(p2741,p2658,p2746,p2747);
HA ha479(p2660,p2743,p2748,p2749);
HA ha480(p2745,p2662,p2750,p2751);
HA ha481(p2664,p2747,p2752,p2753);
HA ha482(p2749,p2666,p2754,p2755);
HA ha483(p2668,p2751,p2756,p2757);
HA ha484(p2753,p2672,p2758,p2759);
HA ha485(p2755,p2757,p2760,p2761);
HA ha486(p2674,p2759,p2762,p2763);
HA ha487(p2761,p2670,p2764,p2765);
HA ha488(p2676,p2678,p2766,p2767);
HA ha489(p2763,p2680,p2768,p2769);
HA ha490(p2682,p2765,p2770,p2771);
HA ha491(p2767,p2684,p2772,p2773);
HA ha492(p2686,p2769,p2774,p2775);
HA ha493(p2771,p2688,p2776,p2777);
HA ha494(p2690,p2773,p2778,p2779);
HA ha495(p2775,p2692,p2780,p2781);
HA ha496(p2694,p2777,p2782,p2783);
HA ha497(p2779,p2696,p2784,p2785);
HA ha498(p2698,p2781,p2786,p2787);
HA ha499(p2783,p2700,p2788,p2789);
HA ha500(p2785,p2787,p2790,p2791);
HA ha501(p2702,p2789,p2792,p2793);
HA ha502(p2791,p2704,p2794,p2795);
HA ha503(ip_31_31,p2706,p2796,p2797);
HA ha504(p2708,p2797,p2798,p2799);
HA ha505(p2710,p2799,p2800,p2801);
FA fa895(p2712,p2714,p2801,p2802,p2803);
HA ha506(p2716,p2718,p2804,p2805);
HA ha507(p2803,p2805,p2806,p2807);
HA ha508(p2722,p2807,p2808,p2809);
HA ha509(p2720,p2724,p2810,p2811);
HA ha510(p2726,p2809,p2812,p2813);
HA ha511(p2728,p2730,p2814,p2815);
HA ha512(p2732,p2811,p2816,p2817);
HA ha513(p2813,p2734,p2818,p2819);
HA ha514(p2736,p2815,p2820,p2821);
HA ha515(p2817,p2740,p2822,p2823);
HA ha516(p2819,p2821,p2824,p2825);
HA ha517(p2738,p2742,p2826,p2827);
HA ha518(p2744,p2823,p2828,p2829);
HA ha519(p2825,p2746,p2830,p2831);
HA ha520(p2748,p2827,p2832,p2833);
HA ha521(p2829,p2750,p2834,p2835);
HA ha522(p2752,p2831,p2836,p2837);
HA ha523(p2833,p2754,p2838,p2839);
HA ha524(p2756,p2835,p2840,p2841);
HA ha525(p2837,p2758,p2842,p2843);
HA ha526(p2760,p2839,p2844,p2845);
HA ha527(p2841,p2762,p2846,p2847);
HA ha528(p2843,p2845,p2848,p2849);
HA ha529(p2764,p2766,p2850,p2851);
HA ha530(p2847,p2849,p2852,p2853);
HA ha531(p2768,p2770,p2854,p2855);
HA ha532(p2851,p2853,p2856,p2857);
HA ha533(p2772,p2774,p2858,p2859);
FA fa896(p2855,p2857,p2776,p2860,p2861);
HA ha534(p2778,p2859,p2862,p2863);
HA ha535(p2780,p2782,p2864,p2865);
HA ha536(p2861,p2863,p2866,p2867);
HA ha537(p2784,p2786,p2868,p2869);
HA ha538(p2865,p2867,p2870,p2871);
HA ha539(p2788,p2790,p2872,p2873);
HA ha540(p2869,p2871,p2874,p2875);
HA ha541(p2792,p2873,p2876,p2877);
HA ha542(p2875,p2794,p2878,p2879);
wire [63:0] a,b;
wire [63:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p5;
assign b[3] = 1'b0;
assign a[4] = p11;
assign b[4] = 1'b0;
assign a[5] = p19;
assign b[5] = 1'b0;
assign a[6] = p29;
assign b[6] = 1'b0;
assign a[7] = p41;
assign b[7] = 1'b0;
assign a[8] = p55;
assign b[8] = 1'b0;
assign a[9] = p71;
assign b[9] = 1'b0;
assign a[10] = p89;
assign b[10] = 1'b0;
assign a[11] = p109;
assign b[11] = 1'b0;
assign a[12] = p131;
assign b[12] = 1'b0;
assign a[13] = p155;
assign b[13] = 1'b0;
assign a[14] = p181;
assign b[14] = 1'b0;
assign a[15] = p209;
assign b[15] = 1'b0;
assign a[16] = p239;
assign b[16] = 1'b0;
assign a[17] = p271;
assign b[17] = 1'b0;
assign a[18] = p305;
assign b[18] = 1'b0;
assign a[19] = p341;
assign b[19] = 1'b0;
assign a[20] = p379;
assign b[20] = 1'b0;
assign a[21] = p419;
assign b[21] = 1'b0;
assign a[22] = p461;
assign b[22] = 1'b0;
assign a[23] = p505;
assign b[23] = 1'b0;
assign a[24] = p551;
assign b[24] = 1'b0;
assign a[25] = p599;
assign b[25] = 1'b0;
assign a[26] = p649;
assign b[26] = 1'b0;
assign a[27] = p701;
assign b[27] = 1'b0;
assign a[28] = p755;
assign b[28] = 1'b0;
assign a[29] = p811;
assign b[29] = p754;
assign a[30] = p869;
assign b[30] = 1'b0;
assign a[31] = p929;
assign b[31] = 1'b0;
assign a[32] = p989;
assign b[32] = 1'b0;
assign a[33] = p1049;
assign b[33] = 1'b0;
assign a[34] = p1107;
assign b[34] = 1'b0;
assign a[35] = p1163;
assign b[35] = 1'b0;
assign a[36] = p1217;
assign b[36] = 1'b0;
assign a[37] = p1269;
assign b[37] = 1'b0;
assign a[38] = p1321;
assign b[38] = 1'b0;
assign a[39] = p1369;
assign b[39] = p1320;
assign a[40] = p1415;
assign b[40] = p1368;
assign a[41] = p1463;
assign b[41] = 1'b0;
assign a[42] = p1511;
assign b[42] = 1'b0;
assign a[43] = p1557;
assign b[43] = 1'b0;
assign a[44] = p1599;
assign b[44] = p1556;
assign a[45] = p1641;
assign b[45] = p1598;
assign a[46] = p1683;
assign b[46] = p1640;
assign a[47] = p1729;
assign b[47] = 1'b0;
assign a[48] = p1773;
assign b[48] = p1728;
assign a[49] = p1825;
assign b[49] = p1772;
assign a[50] = p1881;
assign b[50] = p1824;
assign a[51] = p1943;
assign b[51] = p1880;
assign a[52] = p1942;
assign b[52] = p2005;
assign a[53] = p2004;
assign b[53] = p2077;
assign a[54] = p2151;
assign b[54] = p2153;
assign a[55] = p2239;
assign b[55] = p2241;
assign a[56] = p2327;
assign b[56] = p2329;
assign a[57] = p2326;
assign b[57] = p2423;
assign a[58] = p2515;
assign b[58] = p2517;
assign a[59] = p2609;
assign b[59] = p2611;
assign a[60] = p2703;
assign b[60] = p2705;
assign a[61] = p2793;
assign b[61] = p2795;
assign a[62] = p2877;
assign b[62] = p2879;
assign a[63] = p2796;
assign b[63] = p2798;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[63] = s[63] & p2800 & p2804 & p2802 & p2806 & p2808 & p2810 & p2812 & p2814 & p2816 & p2818 & p2820 & p2822 & p2824 & p2826 & p2828 & p2830 & p2832 & p2834 & p2836 & p2838 & p2840 & p2842 & p2844 & p2846 & p2848 & p2850 & p2852 & p2854 & p2856 & p2858 & p2862 & p2860 & p2864 & p2866 & p2868 & p2870 & p2872 & p2874 & p2876 & p2878;
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
assign o[31] = s[31];
assign o[32] = s[32];
assign o[33] = s[33];
assign o[34] = s[34];
assign o[35] = s[35];
assign o[36] = s[36];
assign o[37] = s[37];
assign o[38] = s[38];
assign o[39] = s[39];
assign o[40] = s[40];
assign o[41] = s[41];
assign o[42] = s[42];
assign o[43] = s[43];
assign o[44] = s[44];
assign o[45] = s[45];
assign o[46] = s[46];
assign o[47] = s[47];
assign o[48] = s[48];
assign o[49] = s[49];
assign o[50] = s[50];
assign o[51] = s[51];
assign o[52] = s[52];
assign o[53] = s[53];
assign o[54] = s[54];
assign o[55] = s[55];
assign o[56] = s[56];
assign o[57] = s[57];
assign o[58] = s[58];
assign o[59] = s[59];
assign o[60] = s[60];
assign o[61] = s[61];
assign o[62] = s[62];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 
module adder(a,b,s);
input [63:0] a,b;
output [63:0] s;
wire g9_8,p42_42,c24,g31_31,g3_3,g24_24,c0,p47_47,g8_8,p56_56,g63_56,g63_62,p50_50,p47_44,g7_4,p2_2,g25_25,p53_52,c59,p62_62,p51_51,g11_0,g15_15,c20,c63,c56,g59_59,g1_1,p7_4,p30_30,p41_41,g49_0,c41,g0_0,g53_52,g37_36,g23_16,p47_46,p5_5,g23_23,p23_16,c37,g39_39,g51_0,c60,g45_0,g28_28,p11_8,g5_0,p15_15,g43_0,p0_0,g33_33,g39_36,g27_27,p10_10,g10_10,g63_48,g55_0,c36,p59_56,g61_61,g47_32,g56_56,p54_54,g9_0,p6_6,p27_27,g50_50,g61_0,p36_36,c9,p14_14,g58_58,p63_62,p4_4,p55_54,p31_31,g59_58,p13_12,g53_0,p37_37,g2_2,p45_44,g26_26,c35,c10,g41_0,g7_7,g62_62,p25_24,p28_28,g17_16,p26_26,g25_24,p33_33,p29_29,g11_11,p59_58,g32_32,p13_13,c58,p31_28,p55_48,g63_32,p11_11,p45_45,p21_21,g19_19,g37_0,c22,c39,g63_63,g54_54,g43_43,g59_56,g5_4,c1,g25_0,p38_38,p11_10,p48_48,g33_0,p44_44,p31_30,p21_20,p49_48,g18_18,c61,g43_40,g57_0,g13_0,g3_0,p57_56,g6_6,c11,g31_16,g38_38,p43_43,g27_0,p51_50,p43_42,p34_34,p22_22,c4,p25_25,g19_0,p7_7,g21_20,c28,c14,c19,c29,g27_24,g31_30,c34,g29_28,g51_50,c53,p23_23,c13,p32_32,c57,g4_4,p15_14,g63_60,p31_24,g14_14,g13_12,g7_0,g20_20,p19_18,p52_52,p12_12,c16,p39_36,c55,p24_24,c38,p16_16,p63_32,p35_34,p47_40,c3,g15_14,g39_0,g22_22,p47_32,c23,p60_60,p15_12,g44_44,g39_38,g7_6,c54,p53_53,g34_34,c8,g3_2,g35_34,c47,c33,c25,c26,p39_39,g43_42,c49,g15_8,g52_52,g47_47,p61_61,g57_57,g37_37,c18,g41_41,p57_57,p17_17,g41_40,g17_17,p1_1,g17_0,c7,c48,c50,g19_16,g61_60,c52,g36_36,p33_32,g15_0,c44,g31_28,g42_42,c21,g11_10,g47_44,c42,c5,c46,g30_30,p7_6,c27,g31_24,g21_21,g35_32,g39_32,p39_38,c62,c30,g35_0,g49_48,p23_22,g51_51,p19_19,g29_29,g55_55,g55_54,p20_20,p9_9,p3_2,p63_56,p61_60,p18_18,p59_59,c17,g40_40,g1_0,p19_16,g53_53,c43,p55_55,g46_46,g16_16,g47_46,g47_0,g19_18,c32,p29_28,g55_52,g35_35,g60_60,c12,c40,g59_0,p27_26,p63_48,p43_40,g9_9,g31_0,g23_22,p41_40,p63_63,g23_20,p27_24,p58_58,c6,g23_0,p51_48,g27_26,g51_48,p40_40,g12_12,c51,p5_4,c2,p35_35,g15_12,g48_48,p55_52,p49_49,g29_0,p9_8,p3_3,g45_44,p63_60,g45_45,p46_46,g49_49,g21_0,p39_32,c31,p17_16,g55_48,p37_36,g47_40,c15,p8_8,g57_56,g5_5,p35_32,g11_8,p23_20,c45,p31_16,p15_8,g33_32,g13_13;

assign p0_0 = a[0] ^ b[0];
assign g0_0 = a[0] & b[0];
assign p1_1 = a[1] ^ b[1];
assign g1_1 = a[1] & b[1];
assign p2_2 = a[2] ^ b[2];
assign g2_2 = a[2] & b[2];
assign p3_3 = a[3] ^ b[3];
assign g3_3 = a[3] & b[3];
assign p4_4 = a[4] ^ b[4];
assign g4_4 = a[4] & b[4];
assign p5_5 = a[5] ^ b[5];
assign g5_5 = a[5] & b[5];
assign p6_6 = a[6] ^ b[6];
assign g6_6 = a[6] & b[6];
assign p7_7 = a[7] ^ b[7];
assign g7_7 = a[7] & b[7];
assign p8_8 = a[8] ^ b[8];
assign g8_8 = a[8] & b[8];
assign p9_9 = a[9] ^ b[9];
assign g9_9 = a[9] & b[9];
assign p10_10 = a[10] ^ b[10];
assign g10_10 = a[10] & b[10];
assign p11_11 = a[11] ^ b[11];
assign g11_11 = a[11] & b[11];
assign p12_12 = a[12] ^ b[12];
assign g12_12 = a[12] & b[12];
assign p13_13 = a[13] ^ b[13];
assign g13_13 = a[13] & b[13];
assign p14_14 = a[14] ^ b[14];
assign g14_14 = a[14] & b[14];
assign p15_15 = a[15] ^ b[15];
assign g15_15 = a[15] & b[15];
assign p16_16 = a[16] ^ b[16];
assign g16_16 = a[16] & b[16];
assign p17_17 = a[17] ^ b[17];
assign g17_17 = a[17] & b[17];
assign p18_18 = a[18] ^ b[18];
assign g18_18 = a[18] & b[18];
assign p19_19 = a[19] ^ b[19];
assign g19_19 = a[19] & b[19];
assign p20_20 = a[20] ^ b[20];
assign g20_20 = a[20] & b[20];
assign p21_21 = a[21] ^ b[21];
assign g21_21 = a[21] & b[21];
assign p22_22 = a[22] ^ b[22];
assign g22_22 = a[22] & b[22];
assign p23_23 = a[23] ^ b[23];
assign g23_23 = a[23] & b[23];
assign p24_24 = a[24] ^ b[24];
assign g24_24 = a[24] & b[24];
assign p25_25 = a[25] ^ b[25];
assign g25_25 = a[25] & b[25];
assign p26_26 = a[26] ^ b[26];
assign g26_26 = a[26] & b[26];
assign p27_27 = a[27] ^ b[27];
assign g27_27 = a[27] & b[27];
assign p28_28 = a[28] ^ b[28];
assign g28_28 = a[28] & b[28];
assign p29_29 = a[29] ^ b[29];
assign g29_29 = a[29] & b[29];
assign p30_30 = a[30] ^ b[30];
assign g30_30 = a[30] & b[30];
assign p31_31 = a[31] ^ b[31];
assign g31_31 = a[31] & b[31];
assign p32_32 = a[32] ^ b[32];
assign g32_32 = a[32] & b[32];
assign p33_33 = a[33] ^ b[33];
assign g33_33 = a[33] & b[33];
assign p34_34 = a[34] ^ b[34];
assign g34_34 = a[34] & b[34];
assign p35_35 = a[35] ^ b[35];
assign g35_35 = a[35] & b[35];
assign p36_36 = a[36] ^ b[36];
assign g36_36 = a[36] & b[36];
assign p37_37 = a[37] ^ b[37];
assign g37_37 = a[37] & b[37];
assign p38_38 = a[38] ^ b[38];
assign g38_38 = a[38] & b[38];
assign p39_39 = a[39] ^ b[39];
assign g39_39 = a[39] & b[39];
assign p40_40 = a[40] ^ b[40];
assign g40_40 = a[40] & b[40];
assign p41_41 = a[41] ^ b[41];
assign g41_41 = a[41] & b[41];
assign p42_42 = a[42] ^ b[42];
assign g42_42 = a[42] & b[42];
assign p43_43 = a[43] ^ b[43];
assign g43_43 = a[43] & b[43];
assign p44_44 = a[44] ^ b[44];
assign g44_44 = a[44] & b[44];
assign p45_45 = a[45] ^ b[45];
assign g45_45 = a[45] & b[45];
assign p46_46 = a[46] ^ b[46];
assign g46_46 = a[46] & b[46];
assign p47_47 = a[47] ^ b[47];
assign g47_47 = a[47] & b[47];
assign p48_48 = a[48] ^ b[48];
assign g48_48 = a[48] & b[48];
assign p49_49 = a[49] ^ b[49];
assign g49_49 = a[49] & b[49];
assign p50_50 = a[50] ^ b[50];
assign g50_50 = a[50] & b[50];
assign p51_51 = a[51] ^ b[51];
assign g51_51 = a[51] & b[51];
assign p52_52 = a[52] ^ b[52];
assign g52_52 = a[52] & b[52];
assign p53_53 = a[53] ^ b[53];
assign g53_53 = a[53] & b[53];
assign p54_54 = a[54] ^ b[54];
assign g54_54 = a[54] & b[54];
assign p55_55 = a[55] ^ b[55];
assign g55_55 = a[55] & b[55];
assign p56_56 = a[56] ^ b[56];
assign g56_56 = a[56] & b[56];
assign p57_57 = a[57] ^ b[57];
assign g57_57 = a[57] & b[57];
assign p58_58 = a[58] ^ b[58];
assign g58_58 = a[58] & b[58];
assign p59_59 = a[59] ^ b[59];
assign g59_59 = a[59] & b[59];
assign p60_60 = a[60] ^ b[60];
assign g60_60 = a[60] & b[60];
assign p61_61 = a[61] ^ b[61];
assign g61_61 = a[61] & b[61];
assign p62_62 = a[62] ^ b[62];
assign g62_62 = a[62] & b[62];
assign p63_63 = a[63] ^ b[63];
assign g63_63 = a[63] & b[63];
assign g1_0 = c1;
assign g2_0 = c2;
assign g3_0 = c3;
assign g4_0 = c4;
assign g5_0 = c5;
assign g6_0 = c6;
assign g7_0 = c7;
assign g8_0 = c8;
assign g9_0 = c9;
assign g10_0 = c10;
assign g11_0 = c11;
assign g12_0 = c12;
assign g13_0 = c13;
assign g14_0 = c14;
assign g15_0 = c15;
assign g16_0 = c16;
assign g17_0 = c17;
assign g18_0 = c18;
assign g19_0 = c19;
assign g20_0 = c20;
assign g21_0 = c21;
assign g22_0 = c22;
assign g23_0 = c23;
assign g24_0 = c24;
assign g25_0 = c25;
assign g26_0 = c26;
assign g27_0 = c27;
assign g28_0 = c28;
assign g29_0 = c29;
assign g30_0 = c30;
assign g31_0 = c31;
assign g32_0 = c32;
assign g33_0 = c33;
assign g34_0 = c34;
assign g35_0 = c35;
assign g36_0 = c36;
assign g37_0 = c37;
assign g38_0 = c38;
assign g39_0 = c39;
assign g40_0 = c40;
assign g41_0 = c41;
assign g42_0 = c42;
assign g43_0 = c43;
assign g44_0 = c44;
assign g45_0 = c45;
assign g46_0 = c46;
assign g47_0 = c47;
assign g48_0 = c48;
assign g49_0 = c49;
assign g50_0 = c50;
assign g51_0 = c51;
assign g52_0 = c52;
assign g53_0 = c53;
assign g54_0 = c54;
assign g55_0 = c55;
assign g56_0 = c56;
assign g57_0 = c57;
assign g58_0 = c58;
assign g59_0 = c59;
assign g60_0 = c60;
assign g61_0 = c61;
assign g62_0 = c62;
assign g63_0 = c63;
BLACK black63_62(g63_63, p63_63, g62_62, p62_62, g63_62, p63_62);
BLACK black63_60(g63_62, p63_62, g61_60, p61_60, g63_60, p63_60);
BLACK black63_56(g63_60, p63_60, g59_56, p59_56, g63_56, p63_56);
BLACK black63_48(g63_56, p63_56, g55_48, p55_48, g63_48, p63_48);
BLACK black63_32(g63_48, p63_48, g47_32, p47_32, g63_32, p63_32);
GREY grey63(g63_32, p63_32, g31_0, c63);
GREY grey62(g62_62, p62_62, g61_0, c62);
BLACK black61_60(g61_61, p61_61, g60_60, p60_60, g61_60, p61_60);
GREY grey61(g61_60, p61_60, g59_0, c61);
GREY grey60(g60_60, p60_60, g59_0, c60);
BLACK black59_58(g59_59, p59_59, g58_58, p58_58, g59_58, p59_58);
BLACK black59_56(g59_58, p59_58, g57_56, p57_56, g59_56, p59_56);
GREY grey59(g59_56, p59_56, g55_0, c59);
GREY grey58(g58_58, p58_58, g57_0, c58);
BLACK black57_56(g57_57, p57_57, g56_56, p56_56, g57_56, p57_56);
GREY grey57(g57_56, p57_56, g55_0, c57);
GREY grey56(g56_56, p56_56, g55_0, c56);
BLACK black55_54(g55_55, p55_55, g54_54, p54_54, g55_54, p55_54);
BLACK black55_52(g55_54, p55_54, g53_52, p53_52, g55_52, p55_52);
BLACK black55_48(g55_52, p55_52, g51_48, p51_48, g55_48, p55_48);
GREY grey55(g55_48, p55_48, g47_0, c55);
GREY grey54(g54_54, p54_54, g53_0, c54);
BLACK black53_52(g53_53, p53_53, g52_52, p52_52, g53_52, p53_52);
GREY grey53(g53_52, p53_52, g51_0, c53);
GREY grey52(g52_52, p52_52, g51_0, c52);
BLACK black51_50(g51_51, p51_51, g50_50, p50_50, g51_50, p51_50);
BLACK black51_48(g51_50, p51_50, g49_48, p49_48, g51_48, p51_48);
GREY grey51(g51_48, p51_48, g47_0, c51);
GREY grey50(g50_50, p50_50, g49_0, c50);
BLACK black49_48(g49_49, p49_49, g48_48, p48_48, g49_48, p49_48);
GREY grey49(g49_48, p49_48, g47_0, c49);
GREY grey48(g48_48, p48_48, g47_0, c48);
BLACK black47_46(g47_47, p47_47, g46_46, p46_46, g47_46, p47_46);
BLACK black47_44(g47_46, p47_46, g45_44, p45_44, g47_44, p47_44);
BLACK black47_40(g47_44, p47_44, g43_40, p43_40, g47_40, p47_40);
BLACK black47_32(g47_40, p47_40, g39_32, p39_32, g47_32, p47_32);
GREY grey47(g47_32, p47_32, g31_0, c47);
GREY grey46(g46_46, p46_46, g45_0, c46);
BLACK black45_44(g45_45, p45_45, g44_44, p44_44, g45_44, p45_44);
GREY grey45(g45_44, p45_44, g43_0, c45);
GREY grey44(g44_44, p44_44, g43_0, c44);
BLACK black43_42(g43_43, p43_43, g42_42, p42_42, g43_42, p43_42);
BLACK black43_40(g43_42, p43_42, g41_40, p41_40, g43_40, p43_40);
GREY grey43(g43_40, p43_40, g39_0, c43);
GREY grey42(g42_42, p42_42, g41_0, c42);
BLACK black41_40(g41_41, p41_41, g40_40, p40_40, g41_40, p41_40);
GREY grey41(g41_40, p41_40, g39_0, c41);
GREY grey40(g40_40, p40_40, g39_0, c40);
BLACK black39_38(g39_39, p39_39, g38_38, p38_38, g39_38, p39_38);
BLACK black39_36(g39_38, p39_38, g37_36, p37_36, g39_36, p39_36);
BLACK black39_32(g39_36, p39_36, g35_32, p35_32, g39_32, p39_32);
GREY grey39(g39_32, p39_32, g31_0, c39);
GREY grey38(g38_38, p38_38, g37_0, c38);
BLACK black37_36(g37_37, p37_37, g36_36, p36_36, g37_36, p37_36);
GREY grey37(g37_36, p37_36, g35_0, c37);
GREY grey36(g36_36, p36_36, g35_0, c36);
BLACK black35_34(g35_35, p35_35, g34_34, p34_34, g35_34, p35_34);
BLACK black35_32(g35_34, p35_34, g33_32, p33_32, g35_32, p35_32);
GREY grey35(g35_32, p35_32, g31_0, c35);
GREY grey34(g34_34, p34_34, g33_0, c34);
BLACK black33_32(g33_33, p33_33, g32_32, p32_32, g33_32, p33_32);
GREY grey33(g33_32, p33_32, g31_0, c33);
GREY grey32(g32_32, p32_32, g31_0, c32);
BLACK black31_30(g31_31, p31_31, g30_30, p30_30, g31_30, p31_30);
BLACK black31_28(g31_30, p31_30, g29_28, p29_28, g31_28, p31_28);
BLACK black31_24(g31_28, p31_28, g27_24, p27_24, g31_24, p31_24);
BLACK black31_16(g31_24, p31_24, g23_16, p23_16, g31_16, p31_16);
GREY grey31(g31_16, p31_16, g15_0, c31);
GREY grey30(g30_30, p30_30, g29_0, c30);
BLACK black29_28(g29_29, p29_29, g28_28, p28_28, g29_28, p29_28);
GREY grey29(g29_28, p29_28, g27_0, c29);
GREY grey28(g28_28, p28_28, g27_0, c28);
BLACK black27_26(g27_27, p27_27, g26_26, p26_26, g27_26, p27_26);
BLACK black27_24(g27_26, p27_26, g25_24, p25_24, g27_24, p27_24);
GREY grey27(g27_24, p27_24, g23_0, c27);
GREY grey26(g26_26, p26_26, g25_0, c26);
BLACK black25_24(g25_25, p25_25, g24_24, p24_24, g25_24, p25_24);
GREY grey25(g25_24, p25_24, g23_0, c25);
GREY grey24(g24_24, p24_24, g23_0, c24);
BLACK black23_22(g23_23, p23_23, g22_22, p22_22, g23_22, p23_22);
BLACK black23_20(g23_22, p23_22, g21_20, p21_20, g23_20, p23_20);
BLACK black23_16(g23_20, p23_20, g19_16, p19_16, g23_16, p23_16);
GREY grey23(g23_16, p23_16, g15_0, c23);
GREY grey22(g22_22, p22_22, g21_0, c22);
BLACK black21_20(g21_21, p21_21, g20_20, p20_20, g21_20, p21_20);
GREY grey21(g21_20, p21_20, g19_0, c21);
GREY grey20(g20_20, p20_20, g19_0, c20);
BLACK black19_18(g19_19, p19_19, g18_18, p18_18, g19_18, p19_18);
BLACK black19_16(g19_18, p19_18, g17_16, p17_16, g19_16, p19_16);
GREY grey19(g19_16, p19_16, g15_0, c19);
GREY grey18(g18_18, p18_18, g17_0, c18);
BLACK black17_16(g17_17, p17_17, g16_16, p16_16, g17_16, p17_16);
GREY grey17(g17_16, p17_16, g15_0, c17);
GREY grey16(g16_16, p16_16, g15_0, c16);
BLACK black15_14(g15_15, p15_15, g14_14, p14_14, g15_14, p15_14);
BLACK black15_12(g15_14, p15_14, g13_12, p13_12, g15_12, p15_12);
BLACK black15_8(g15_12, p15_12, g11_8, p11_8, g15_8, p15_8);
GREY grey15(g15_8, p15_8, g7_0, c15);
GREY grey14(g14_14, p14_14, g13_0, c14);
BLACK black13_12(g13_13, p13_13, g12_12, p12_12, g13_12, p13_12);
GREY grey13(g13_12, p13_12, g11_0, c13);
GREY grey12(g12_12, p12_12, g11_0, c12);
BLACK black11_10(g11_11, p11_11, g10_10, p10_10, g11_10, p11_10);
BLACK black11_8(g11_10, p11_10, g9_8, p9_8, g11_8, p11_8);
GREY grey11(g11_8, p11_8, g7_0, c11);
GREY grey10(g10_10, p10_10, g9_0, c10);
BLACK black9_8(g9_9, p9_9, g8_8, p8_8, g9_8, p9_8);
GREY grey9(g9_8, p9_8, g7_0, c9);
GREY grey8(g8_8, p8_8, g7_0, c8);
BLACK black7_6(g7_7, p7_7, g6_6, p6_6, g7_6, p7_6);
BLACK black7_4(g7_6, p7_6, g5_4, p5_4, g7_4, p7_4);
GREY grey7(g7_4, p7_4, g3_0, c7);
GREY grey6(g6_6, p6_6, g5_0, c6);
BLACK black5_4(g5_5, p5_5, g4_4, p4_4, g5_4, p5_4);
GREY grey5(g5_4, p5_4, g3_0, c5);
GREY grey4(g4_4, p4_4, g3_0, c4);
BLACK black3_2(g3_3, p3_3, g2_2, p2_2, g3_2, p3_2);
GREY grey3(g3_2, p3_2, g1_0, c3);
GREY grey2(g2_2, p2_2, g1_0, c2);
GREY grey1(g1_1, p1_1, g0_0, c1);
assign s[0] = a[0] ^ b[0];
assign c0 = g0_0;
assign s[1] = p1_1 ^ c0;
assign s[2] = p2_2 ^ c1;
assign s[3] = p3_3 ^ c2;
assign s[4] = p4_4 ^ c3;
assign s[5] = p5_5 ^ c4;
assign s[6] = p6_6 ^ c5;
assign s[7] = p7_7 ^ c6;
assign s[8] = p8_8 ^ c7;
assign s[9] = p9_9 ^ c8;
assign s[10] = p10_10 ^ c9;
assign s[11] = p11_11 ^ c10;
assign s[12] = p12_12 ^ c11;
assign s[13] = p13_13 ^ c12;
assign s[14] = p14_14 ^ c13;
assign s[15] = p15_15 ^ c14;
assign s[16] = p16_16 ^ c15;
assign s[17] = p17_17 ^ c16;
assign s[18] = p18_18 ^ c17;
assign s[19] = p19_19 ^ c18;
assign s[20] = p20_20 ^ c19;
assign s[21] = p21_21 ^ c20;
assign s[22] = p22_22 ^ c21;
assign s[23] = p23_23 ^ c22;
assign s[24] = p24_24 ^ c23;
assign s[25] = p25_25 ^ c24;
assign s[26] = p26_26 ^ c25;
assign s[27] = p27_27 ^ c26;
assign s[28] = p28_28 ^ c27;
assign s[29] = p29_29 ^ c28;
assign s[30] = p30_30 ^ c29;
assign s[31] = p31_31 ^ c30;
assign s[32] = p32_32 ^ c31;
assign s[33] = p33_33 ^ c32;
assign s[34] = p34_34 ^ c33;
assign s[35] = p35_35 ^ c34;
assign s[36] = p36_36 ^ c35;
assign s[37] = p37_37 ^ c36;
assign s[38] = p38_38 ^ c37;
assign s[39] = p39_39 ^ c38;
assign s[40] = p40_40 ^ c39;
assign s[41] = p41_41 ^ c40;
assign s[42] = p42_42 ^ c41;
assign s[43] = p43_43 ^ c42;
assign s[44] = p44_44 ^ c43;
assign s[45] = p45_45 ^ c44;
assign s[46] = p46_46 ^ c45;
assign s[47] = p47_47 ^ c46;
assign s[48] = p48_48 ^ c47;
assign s[49] = p49_49 ^ c48;
assign s[50] = p50_50 ^ c49;
assign s[51] = p51_51 ^ c50;
assign s[52] = p52_52 ^ c51;
assign s[53] = p53_53 ^ c52;
assign s[54] = p54_54 ^ c53;
assign s[55] = p55_55 ^ c54;
assign s[56] = p56_56 ^ c55;
assign s[57] = p57_57 ^ c56;
assign s[58] = p58_58 ^ c57;
assign s[59] = p59_59 ^ c58;
assign s[60] = p60_60 ^ c59;
assign s[61] = p61_61 ^ c60;
assign s[62] = p62_62 ^ c61;
assign s[63] = p63_63 ^ c62;
endmodule

module GREY(gik, pik, gkj, gij);
input gik, pik, gkj;
output gij;
assign gij = gik | (pik & gkj);
endmodule

module BLACK(gik, pik, gkj, pkj, gij, pij);
input gik, pik, gkj, pkj;
output gij, pij;
assign pij = pik & pkj;
assign gij = gik | (pik & gkj);
endmodule

