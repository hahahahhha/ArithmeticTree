// 1 2 1 2 2 2 2 1 2 1 2 2 2 2 2 2 2 2 2 1 2 1 2 3 

module main(x,y,o);
input [11:0] x,y;
output [23:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_1_0,x[1],y[0]);
and and13(ip_1_1,x[1],y[1]);
and and14(ip_1_2,x[1],y[2]);
and and15(ip_1_3,x[1],y[3]);
and and16(ip_1_4,x[1],y[4]);
and and17(ip_1_5,x[1],y[5]);
and and18(ip_1_6,x[1],y[6]);
and and19(ip_1_7,x[1],y[7]);
and and20(ip_1_8,x[1],y[8]);
and and21(ip_1_9,x[1],y[9]);
and and22(ip_1_10,x[1],y[10]);
and and23(ip_1_11,x[1],y[11]);
and and24(ip_2_0,x[2],y[0]);
and and25(ip_2_1,x[2],y[1]);
and and26(ip_2_2,x[2],y[2]);
and and27(ip_2_3,x[2],y[3]);
and and28(ip_2_4,x[2],y[4]);
and and29(ip_2_5,x[2],y[5]);
and and30(ip_2_6,x[2],y[6]);
and and31(ip_2_7,x[2],y[7]);
and and32(ip_2_8,x[2],y[8]);
and and33(ip_2_9,x[2],y[9]);
and and34(ip_2_10,x[2],y[10]);
and and35(ip_2_11,x[2],y[11]);
and and36(ip_3_0,x[3],y[0]);
and and37(ip_3_1,x[3],y[1]);
and and38(ip_3_2,x[3],y[2]);
and and39(ip_3_3,x[3],y[3]);
and and40(ip_3_4,x[3],y[4]);
and and41(ip_3_5,x[3],y[5]);
and and42(ip_3_6,x[3],y[6]);
and and43(ip_3_7,x[3],y[7]);
and and44(ip_3_8,x[3],y[8]);
and and45(ip_3_9,x[3],y[9]);
and and46(ip_3_10,x[3],y[10]);
and and47(ip_3_11,x[3],y[11]);
and and48(ip_4_0,x[4],y[0]);
and and49(ip_4_1,x[4],y[1]);
and and50(ip_4_2,x[4],y[2]);
and and51(ip_4_3,x[4],y[3]);
and and52(ip_4_4,x[4],y[4]);
and and53(ip_4_5,x[4],y[5]);
and and54(ip_4_6,x[4],y[6]);
and and55(ip_4_7,x[4],y[7]);
and and56(ip_4_8,x[4],y[8]);
and and57(ip_4_9,x[4],y[9]);
and and58(ip_4_10,x[4],y[10]);
and and59(ip_4_11,x[4],y[11]);
and and60(ip_5_0,x[5],y[0]);
and and61(ip_5_1,x[5],y[1]);
and and62(ip_5_2,x[5],y[2]);
and and63(ip_5_3,x[5],y[3]);
and and64(ip_5_4,x[5],y[4]);
and and65(ip_5_5,x[5],y[5]);
and and66(ip_5_6,x[5],y[6]);
and and67(ip_5_7,x[5],y[7]);
and and68(ip_5_8,x[5],y[8]);
and and69(ip_5_9,x[5],y[9]);
and and70(ip_5_10,x[5],y[10]);
and and71(ip_5_11,x[5],y[11]);
and and72(ip_6_0,x[6],y[0]);
and and73(ip_6_1,x[6],y[1]);
and and74(ip_6_2,x[6],y[2]);
and and75(ip_6_3,x[6],y[3]);
and and76(ip_6_4,x[6],y[4]);
and and77(ip_6_5,x[6],y[5]);
and and78(ip_6_6,x[6],y[6]);
and and79(ip_6_7,x[6],y[7]);
and and80(ip_6_8,x[6],y[8]);
and and81(ip_6_9,x[6],y[9]);
and and82(ip_6_10,x[6],y[10]);
and and83(ip_6_11,x[6],y[11]);
and and84(ip_7_0,x[7],y[0]);
and and85(ip_7_1,x[7],y[1]);
and and86(ip_7_2,x[7],y[2]);
and and87(ip_7_3,x[7],y[3]);
and and88(ip_7_4,x[7],y[4]);
and and89(ip_7_5,x[7],y[5]);
and and90(ip_7_6,x[7],y[6]);
and and91(ip_7_7,x[7],y[7]);
and and92(ip_7_8,x[7],y[8]);
and and93(ip_7_9,x[7],y[9]);
and and94(ip_7_10,x[7],y[10]);
and and95(ip_7_11,x[7],y[11]);
and and96(ip_8_0,x[8],y[0]);
and and97(ip_8_1,x[8],y[1]);
and and98(ip_8_2,x[8],y[2]);
and and99(ip_8_3,x[8],y[3]);
and and100(ip_8_4,x[8],y[4]);
and and101(ip_8_5,x[8],y[5]);
and and102(ip_8_6,x[8],y[6]);
and and103(ip_8_7,x[8],y[7]);
and and104(ip_8_8,x[8],y[8]);
and and105(ip_8_9,x[8],y[9]);
and and106(ip_8_10,x[8],y[10]);
and and107(ip_8_11,x[8],y[11]);
and and108(ip_9_0,x[9],y[0]);
and and109(ip_9_1,x[9],y[1]);
and and110(ip_9_2,x[9],y[2]);
and and111(ip_9_3,x[9],y[3]);
and and112(ip_9_4,x[9],y[4]);
and and113(ip_9_5,x[9],y[5]);
and and114(ip_9_6,x[9],y[6]);
and and115(ip_9_7,x[9],y[7]);
and and116(ip_9_8,x[9],y[8]);
and and117(ip_9_9,x[9],y[9]);
and and118(ip_9_10,x[9],y[10]);
and and119(ip_9_11,x[9],y[11]);
and and120(ip_10_0,x[10],y[0]);
and and121(ip_10_1,x[10],y[1]);
and and122(ip_10_2,x[10],y[2]);
and and123(ip_10_3,x[10],y[3]);
and and124(ip_10_4,x[10],y[4]);
and and125(ip_10_5,x[10],y[5]);
and and126(ip_10_6,x[10],y[6]);
and and127(ip_10_7,x[10],y[7]);
and and128(ip_10_8,x[10],y[8]);
and and129(ip_10_9,x[10],y[9]);
and and130(ip_10_10,x[10],y[10]);
and and131(ip_10_11,x[10],y[11]);
and and132(ip_11_0,x[11],y[0]);
and and133(ip_11_1,x[11],y[1]);
and and134(ip_11_2,x[11],y[2]);
and and135(ip_11_3,x[11],y[3]);
and and136(ip_11_4,x[11],y[4]);
and and137(ip_11_5,x[11],y[5]);
and and138(ip_11_6,x[11],y[6]);
and and139(ip_11_7,x[11],y[7]);
and and140(ip_11_8,x[11],y[8]);
and and141(ip_11_9,x[11],y[9]);
and and142(ip_11_10,x[11],y[10]);
and and143(ip_11_11,x[11],y[11]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
HA ha0(ip_0_3,ip_1_2,p2,p3);
FA fa1(ip_2_1,ip_3_0,p3,p4,p5);
FA fa2(ip_0_4,ip_1_3,ip_2_2,p6,p7);
HA ha1(ip_3_1,ip_4_0,p8,p9);
HA ha2(p2,p9,p10,p11);
HA ha3(p11,p7,p12,p13);
HA ha4(ip_0_5,ip_1_4,p14,p15);
FA fa3(ip_2_3,ip_3_2,ip_4_1,p16,p17);
HA ha5(ip_5_0,p15,p18,p19);
FA fa4(p8,p10,p17,p20,p21);
HA ha6(p19,p12,p22,p23);
HA ha7(p6,p21,p24,p25);
HA ha8(ip_0_6,ip_1_5,p26,p27);
HA ha9(ip_2_4,ip_3_3,p28,p29);
HA ha10(ip_4_2,ip_5_1,p30,p31);
FA fa5(ip_6_0,p14,p27,p32,p33);
HA ha11(p29,p31,p34,p35);
FA fa6(p18,p35,p16,p36,p37);
HA ha12(p33,p22,p38,p39);
FA fa7(p37,p20,p24,p40,p41);
FA fa8(ip_0_7,ip_1_6,ip_2_5,p42,p43);
HA ha13(ip_3_4,ip_4_3,p44,p45);
FA fa9(ip_5_2,ip_6_1,ip_7_0,p46,p47);
FA fa10(p26,p28,p30,p48,p49);
HA ha14(p45,p34,p50,p51);
HA ha15(p43,p47,p52,p53);
HA ha16(p49,p51,p54,p55);
HA ha17(p53,p32,p56,p57);
FA fa11(p55,p36,p38,p58,p59);
FA fa12(p57,p59,p40,p60,p61);
HA ha18(ip_0_8,ip_1_7,p62,p63);
HA ha19(ip_2_6,ip_3_5,p64,p65);
HA ha20(ip_4_4,ip_5_3,p66,p67);
HA ha21(ip_6_2,ip_7_1,p68,p69);
FA fa13(ip_8_0,p44,p63,p70,p71);
FA fa14(p65,p67,p69,p72,p73);
HA ha22(p42,p46,p74,p75);
HA ha23(p50,p52,p76,p77);
HA ha24(p71,p73,p78,p79);
HA ha25(p48,p54,p80,p81);
HA ha26(p75,p77,p82,p83);
HA ha27(p79,p56,p84,p85);
HA ha28(p81,p83,p86,p87);
FA fa15(p85,p87,p58,p88,p89);
FA fa16(ip_0_9,ip_1_8,ip_2_7,p90,p91);
FA fa17(ip_3_6,ip_4_5,ip_5_4,p92,p93);
HA ha29(ip_6_3,ip_7_2,p94,p95);
HA ha30(ip_8_1,ip_9_0,p96,p97);
HA ha31(p62,p64,p98,p99);
FA fa18(p66,p68,p95,p100,p101);
FA fa19(p97,p91,p93,p102,p103);
HA ha32(p99,p101,p104,p105);
HA ha33(p103,p105,p106,p107);
FA fa20(p70,p72,p74,p108,p109);
FA fa21(p76,p78,p107,p110,p111);
FA fa22(p80,p82,p109,p112,p113);
HA ha34(p111,p84,p114,p115);
HA ha35(p86,p113,p116,p117);
FA fa23(p115,p117,p88,p118,p119);
HA ha36(ip_0_10,ip_1_9,p120,p121);
FA fa24(ip_2_8,ip_3_7,ip_4_6,p122,p123);
HA ha37(ip_5_5,ip_6_4,p124,p125);
FA fa25(ip_7_3,ip_8_2,ip_9_1,p126,p127);
HA ha38(ip_10_0,p121,p128,p129);
FA fa26(p125,p94,p96,p130,p131);
HA ha39(p123,p127,p132,p133);
HA ha40(p129,p98,p134,p135);
HA ha41(p131,p133,p136,p137);
HA ha42(p135,p90,p138,p139);
FA fa27(p92,p100,p104,p140,p141);
HA ha43(p137,p139,p142,p143);
HA ha44(p102,p106,p144,p145);
HA ha45(p143,p141,p146,p147);
FA fa28(p145,p108,p110,p148,p149);
FA fa29(p114,p147,p112,p150,p151);
FA fa30(p116,p149,p151,p152,p153);
HA ha46(ip_0_11,ip_1_10,p154,p155);
FA fa31(ip_2_9,ip_3_8,ip_4_7,p156,p157);
HA ha47(ip_5_6,ip_6_5,p158,p159);
FA fa32(ip_7_4,ip_8_3,ip_9_2,p160,p161);
FA fa33(ip_10_1,ip_11_0,p120,p162,p163);
HA ha48(p124,p155,p164,p165);
FA fa34(p159,p128,p157,p166,p167);
HA ha49(p161,p163,p168,p169);
FA fa35(p165,p122,p126,p170,p171);
FA fa36(p132,p134,p169,p172,p173);
HA ha50(p130,p136,p174,p175);
HA ha51(p138,p167,p176,p177);
FA fa37(p142,p171,p173,p178,p179);
HA ha52(p175,p177,p180,p181);
FA fa38(p144,p181,p140,p182,p183);
FA fa39(p146,p179,p183,p184,p185);
FA fa40(p185,p148,p150,p186,p187);
FA fa41(ip_1_11,ip_2_10,ip_3_9,p188,p189);
FA fa42(ip_4_8,ip_5_7,ip_6_6,p190,p191);
HA ha53(ip_7_5,ip_8_4,p192,p193);
HA ha54(ip_9_3,ip_10_2,p194,p195);
HA ha55(ip_11_1,p154,p196,p197);
FA fa43(p158,p193,p195,p198,p199);
HA ha56(p164,p189,p200,p201);
FA fa44(p191,p197,p156,p202,p203);
HA ha57(p160,p162,p204,p205);
HA ha58(p168,p199,p206,p207);
FA fa45(p201,p203,p205,p208,p209);
FA fa46(p207,p166,p174,p210,p211);
HA ha59(p176,p170,p212,p213);
FA fa47(p172,p180,p209,p214,p215);
FA fa48(p211,p213,p178,p216,p217);
HA ha60(p215,p182,p218,p219);
FA fa49(p217,p184,p219,p220,p221);
HA ha61(ip_2_11,ip_3_10,p222,p223);
FA fa50(ip_4_9,ip_5_8,ip_6_7,p224,p225);
HA ha62(ip_7_6,ip_8_5,p226,p227);
FA fa51(ip_9_4,ip_10_3,ip_11_2,p228,p229);
HA ha63(p192,p194,p230,p231);
HA ha64(p223,p227,p232,p233);
HA ha65(p196,p225,p234,p235);
FA fa52(p229,p231,p233,p236,p237);
FA fa53(p188,p190,p200,p238,p239);
FA fa54(p235,p198,p204,p240,p241);
FA fa55(p206,p237,p202,p242,p243);
HA ha66(p239,p241,p244,p245);
HA ha67(p243,p208,p246,p247);
HA ha68(p212,p245,p248,p249);
HA ha69(p210,p247,p250,p251);
FA fa56(p249,p214,p251,p252,p253);
FA fa57(p216,p218,p253,p254,p255);
HA ha70(ip_3_11,ip_4_10,p256,p257);
FA fa58(ip_5_9,ip_6_8,ip_7_7,p258,p259);
FA fa59(ip_8_6,ip_9_5,ip_10_4,p260,p261);
FA fa60(ip_11_3,p222,p226,p262,p263);
HA ha71(p257,p230,p264,p265);
FA fa61(p232,p259,p261,p266,p267);
HA ha72(p224,p228,p268,p269);
HA ha73(p234,p263,p270,p271);
HA ha74(p265,p267,p272,p273);
FA fa62(p269,p271,p236,p274,p275);
FA fa63(p273,p238,p275,p276,p277);
FA fa64(p240,p242,p244,p278,p279);
FA fa65(p246,p248,p277,p280,p281);
FA fa66(p250,p279,p281,p282,p283);
HA ha75(p283,p252,p284,p285);
HA ha76(ip_4_11,ip_5_10,p286,p287);
FA fa67(ip_6_9,ip_7_8,ip_8_7,p288,p289);
FA fa68(ip_9_6,ip_10_5,ip_11_4,p290,p291);
FA fa69(p256,p287,p289,p292,p293);
HA ha77(p291,p258,p294,p295);
HA ha78(p260,p264,p296,p297);
FA fa70(p293,p262,p268,p298,p299);
HA ha79(p270,p295,p300,p301);
FA fa71(p297,p266,p272,p302,p303);
FA fa72(p301,p299,p274,p304,p305);
HA ha80(p303,p305,p306,p307);
FA fa73(p276,p307,p278,p308,p309);
FA fa74(p280,p309,p282,p310,p311);
FA fa75(ip_5_11,ip_6_10,ip_7_9,p312,p313);
FA fa76(ip_8_8,ip_9_7,ip_10_6,p314,p315);
FA fa77(ip_11_5,p286,p313,p316,p317);
HA ha81(p315,p288,p318,p319);
FA fa78(p290,p317,p292,p320,p321);
HA ha82(p294,p296,p322,p323);
HA ha83(p319,p300,p324,p325);
HA ha84(p321,p323,p326,p327);
FA fa79(p325,p327,p298,p328,p329);
FA fa80(p302,p329,p304,p330,p331);
HA ha85(p306,p331,p332,p333);
HA ha86(p333,p308,p334,p335);
FA fa81(ip_6_11,ip_7_10,ip_8_9,p336,p337);
FA fa82(ip_9_8,ip_10_7,ip_11_6,p338,p339);
HA ha87(p337,p339,p340,p341);
FA fa83(p312,p314,p341,p342,p343);
FA fa84(p316,p318,p322,p344,p345);
FA fa85(p343,p320,p324,p346,p347);
HA ha88(p326,p345,p348,p349);
HA ha89(p349,p347,p350,p351);
HA ha90(p328,p351,p352,p353);
FA fa86(p353,p330,p332,p354,p355);
FA fa87(ip_7_11,ip_8_10,ip_9_9,p356,p357);
FA fa88(ip_10_8,ip_11_7,p357,p358,p359);
HA ha91(p336,p338,p360,p361);
HA ha92(p340,p359,p362,p363);
HA ha93(p361,p363,p364,p365);
FA fa89(p365,p342,p344,p366,p367);
HA ha94(p348,p367,p368,p369);
FA fa90(p346,p350,p369,p370,p371);
HA ha95(p352,p371,p372,p373);
FA fa91(ip_8_11,ip_9_10,ip_10_9,p374,p375);
HA ha96(ip_11_8,p375,p376,p377);
FA fa92(p356,p377,p358,p378,p379);
FA fa93(p360,p362,p364,p380,p381);
HA ha97(p379,p381,p382,p383);
HA ha98(p383,p366,p384,p385);
HA ha99(p368,p385,p386,p387);
FA fa94(p387,p370,p372,p388,p389);
FA fa95(ip_9_11,ip_10_10,ip_11_9,p390,p391);
HA ha100(p391,p374,p392,p393);
HA ha101(p376,p393,p394,p395);
HA ha102(p395,p378,p396,p397);
HA ha103(p380,p382,p398,p399);
HA ha104(p397,p399,p400,p401);
FA fa96(p401,p384,p386,p402,p403);
FA fa97(ip_10_11,ip_11_10,p390,p404,p405);
FA fa98(p392,p405,p394,p406,p407);
HA ha105(p407,p396,p408,p409);
HA ha106(p398,p409,p410,p411);
FA fa99(p400,p411,p402,p412,p413);
HA ha107(ip_11_11,p404,p414,p415);
FA fa100(p415,p406,p408,p416,p417);
HA ha108(p410,p417,p418,p419);
wire [23:0] a,b;
wire [23:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p5;
assign b[3] = p0;
assign a[4] = p13;
assign b[4] = p4;
assign a[5] = p23;
assign b[5] = p25;
assign a[6] = p39;
assign b[6] = p41;
assign a[7] = p61;
assign b[7] = 1'b0;
assign a[8] = p89;
assign b[8] = p60;
assign a[9] = p119;
assign b[9] = 1'b0;
assign a[10] = p153;
assign b[10] = p118;
assign a[11] = p152;
assign b[11] = p187;
assign a[12] = p221;
assign b[12] = p186;
assign a[13] = p255;
assign b[13] = p220;
assign a[14] = p254;
assign b[14] = p285;
assign a[15] = p284;
assign b[15] = p311;
assign a[16] = p335;
assign b[16] = p310;
assign a[17] = p334;
assign b[17] = p355;
assign a[18] = p373;
assign b[18] = p354;
assign a[19] = p389;
assign b[19] = 1'b0;
assign a[20] = p403;
assign b[20] = p388;
assign a[21] = p413;
assign b[21] = 1'b0;
assign a[22] = p419;
assign b[22] = p412;
assign a[23] = p414;
assign b[23] = p416;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[23] = s[23] & p418;
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [23:0] a,b;
output [23:0] s;
assign s = a+b;
endmodule
