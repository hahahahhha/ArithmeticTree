// 1 2 1 2 2 1 1 2 1 2 2 2 1 2 2 1 

module main(x,y,o);
input [7:0] x,y;
output [15:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_1_0,x[1],y[0]);
and and9(ip_1_1,x[1],y[1]);
and and10(ip_1_2,x[1],y[2]);
and and11(ip_1_3,x[1],y[3]);
and and12(ip_1_4,x[1],y[4]);
and and13(ip_1_5,x[1],y[5]);
and and14(ip_1_6,x[1],y[6]);
and and15(ip_1_7,x[1],y[7]);
and and16(ip_2_0,x[2],y[0]);
and and17(ip_2_1,x[2],y[1]);
and and18(ip_2_2,x[2],y[2]);
and and19(ip_2_3,x[2],y[3]);
and and20(ip_2_4,x[2],y[4]);
and and21(ip_2_5,x[2],y[5]);
and and22(ip_2_6,x[2],y[6]);
and and23(ip_2_7,x[2],y[7]);
and and24(ip_3_0,x[3],y[0]);
and and25(ip_3_1,x[3],y[1]);
and and26(ip_3_2,x[3],y[2]);
and and27(ip_3_3,x[3],y[3]);
and and28(ip_3_4,x[3],y[4]);
and and29(ip_3_5,x[3],y[5]);
and and30(ip_3_6,x[3],y[6]);
and and31(ip_3_7,x[3],y[7]);
and and32(ip_4_0,x[4],y[0]);
and and33(ip_4_1,x[4],y[1]);
and and34(ip_4_2,x[4],y[2]);
and and35(ip_4_3,x[4],y[3]);
and and36(ip_4_4,x[4],y[4]);
and and37(ip_4_5,x[4],y[5]);
and and38(ip_4_6,x[4],y[6]);
and and39(ip_4_7,x[4],y[7]);
and and40(ip_5_0,x[5],y[0]);
and and41(ip_5_1,x[5],y[1]);
and and42(ip_5_2,x[5],y[2]);
and and43(ip_5_3,x[5],y[3]);
and and44(ip_5_4,x[5],y[4]);
and and45(ip_5_5,x[5],y[5]);
and and46(ip_5_6,x[5],y[6]);
and and47(ip_5_7,x[5],y[7]);
and and48(ip_6_0,x[6],y[0]);
and and49(ip_6_1,x[6],y[1]);
and and50(ip_6_2,x[6],y[2]);
and and51(ip_6_3,x[6],y[3]);
and and52(ip_6_4,x[6],y[4]);
and and53(ip_6_5,x[6],y[5]);
and and54(ip_6_6,x[6],y[6]);
and and55(ip_6_7,x[6],y[7]);
and and56(ip_7_0,x[7],y[0]);
and and57(ip_7_1,x[7],y[1]);
and and58(ip_7_2,x[7],y[2]);
and and59(ip_7_3,x[7],y[3]);
and and60(ip_7_4,x[7],y[4]);
and and61(ip_7_5,x[7],y[5]);
and and62(ip_7_6,x[7],y[6]);
and and63(ip_7_7,x[7],y[7]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
HA ha0(ip_3_0,p3,p4,p5);
FA fa2(ip_0_4,ip_1_3,ip_2_2,p6,p7);
HA ha1(ip_3_1,ip_4_0,p8,p9);
FA fa3(p9,p7,p2,p10,p11);
HA ha2(ip_0_5,ip_1_4,p12,p13);
FA fa4(ip_2_3,ip_3_2,ip_4_1,p14,p15);
HA ha3(ip_5_0,p13,p16,p17);
HA ha4(p8,p15,p18,p19);
HA ha5(p17,p19,p20,p21);
FA fa5(p6,p21,p10,p22,p23);
FA fa6(ip_0_6,ip_1_5,ip_2_4,p24,p25);
FA fa7(ip_3_3,ip_4_2,ip_5_1,p26,p27);
FA fa8(ip_6_0,p12,p16,p28,p29);
HA ha6(p25,p27,p30,p31);
HA ha7(p14,p18,p32,p33);
HA ha8(p29,p31,p34,p35);
HA ha9(p20,p33,p36,p37);
FA fa9(p35,p37,p22,p38,p39);
FA fa10(ip_0_7,ip_1_6,ip_2_5,p40,p41);
HA ha10(ip_3_4,ip_4_3,p42,p43);
FA fa11(ip_5_2,ip_6_1,ip_7_0,p44,p45);
FA fa12(p43,p41,p45,p46,p47);
FA fa13(p24,p26,p30,p48,p49);
HA ha11(p28,p32,p50,p51);
FA fa14(p34,p47,p36,p52,p53);
HA ha12(p49,p51,p54,p55);
HA ha13(p53,p55,p56,p57);
HA ha14(ip_1_7,ip_2_6,p58,p59);
FA fa15(ip_3_5,ip_4_4,ip_5_3,p60,p61);
FA fa16(ip_6_2,ip_7_1,p42,p62,p63);
FA fa17(p59,p61,p63,p64,p65);
FA fa18(p40,p44,p65,p66,p67);
FA fa19(p46,p50,p67,p68,p69);
HA ha15(p48,p54,p70,p71);
HA ha16(p52,p56,p72,p73);
FA fa20(p69,p71,p73,p74,p75);
FA fa21(ip_2_7,ip_3_6,ip_4_5,p76,p77);
FA fa22(ip_5_4,ip_6_3,ip_7_2,p78,p79);
HA ha17(p58,p77,p80,p81);
HA ha18(p79,p60,p82,p83);
FA fa23(p62,p81,p83,p84,p85);
HA ha19(p64,p85,p86,p87);
FA fa24(p66,p87,p70,p88,p89);
FA fa25(p68,p72,p89,p90,p91);
HA ha20(ip_3_7,ip_4_6,p92,p93);
FA fa26(ip_5_5,ip_6_4,ip_7_3,p94,p95);
FA fa27(p93,p95,p76,p96,p97);
FA fa28(p78,p80,p82,p98,p99);
FA fa29(p97,p99,p84,p100,p101);
FA fa30(p86,p101,p88,p102,p103);
HA ha21(ip_4_7,ip_5_6,p104,p105);
FA fa31(ip_6_5,ip_7_4,p105,p106,p107);
HA ha22(p92,p107,p108,p109);
HA ha23(p109,p94,p110,p111);
HA ha24(p111,p96,p112,p113);
FA fa32(p113,p98,p100,p114,p115);
FA fa33(ip_5_7,ip_6_6,ip_7_5,p116,p117);
HA ha25(p104,p117,p118,p119);
HA ha26(p106,p108,p120,p121);
FA fa34(p119,p110,p121,p122,p123);
FA fa35(p112,p123,p114,p124,p125);
HA ha27(ip_6_7,ip_7_6,p126,p127);
FA fa36(p127,p116,p118,p128,p129);
FA fa37(p120,p129,p122,p130,p131);
FA fa38(ip_7_7,p126,p128,p132,p133);
wire [15:0] a,b;
wire [15:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p0;
assign b[3] = p5;
assign a[4] = p4;
assign b[4] = p11;
assign a[5] = p23;
assign b[5] = 1'b0;
assign a[6] = p39;
assign b[6] = 1'b0;
assign a[7] = p57;
assign b[7] = p38;
assign a[8] = p75;
assign b[8] = 1'b0;
assign a[9] = p74;
assign b[9] = p91;
assign a[10] = p103;
assign b[10] = p90;
assign a[11] = p115;
assign b[11] = p102;
assign a[12] = p125;
assign b[12] = 1'b0;
assign a[13] = p131;
assign b[13] = p124;
assign a[14] = p133;
assign b[14] = p130;
assign a[15] = p132;
assign b[15] = 1'b0;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[15] = s[15];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [15:0] a,b;
output [15:0] s;
assign s = a+b;
endmodule
