// 1 2 2 2 2 2 2 2 2 1 2 2 2 1 2 1 2 2 2 2 2 2 2 2 2 1 2 2 2 1 1 11 

module main(x,y,o);
input [15:0] x,y;
output [31:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149,p1150,p1151,p1152,p1153,p1154,p1155,p1156,p1157,p1158,p1159,p1160,p1161,p1162,p1163,p1164,p1165,p1166,p1167,p1168,p1169,p1170,p1171,p1172,p1173,p1174,p1175,p1176,p1177,p1178,p1179,p1180,p1181,p1182,p1183,p1184,p1185,p1186,p1187,p1188,p1189,p1190,p1191,p1192,p1193,p1194,p1195,p1196,p1197,p1198,p1199,p1200,p1201,p1202,p1203,p1204,p1205,p1206,p1207,p1208,p1209,p1210,p1211,p1212,p1213,p1214,p1215,p1216,p1217,p1218,p1219,p1220,p1221,p1222,p1223,p1224,p1225,p1226,p1227,p1228,p1229,p1230,p1231,p1232,p1233,p1234,p1235,p1236,p1237,p1238,p1239,p1240,p1241,p1242,p1243,p1244,p1245,p1246,p1247,p1248,p1249,p1250,p1251,p1252,p1253,p1254,p1255,p1256,p1257,p1258,p1259,p1260,p1261,p1262,p1263,p1264,p1265,p1266,p1267,p1268,p1269,p1270,p1271,p1272,p1273,p1274,p1275,p1276,p1277,p1278,p1279,p1280,p1281,p1282,p1283,p1284,p1285,p1286,p1287,p1288,p1289,p1290,p1291,p1292,p1293,p1294,p1295,p1296,p1297,p1298,p1299,p1300,p1301,p1302,p1303,p1304,p1305,p1306,p1307,p1308,p1309,p1310,p1311,p1312,p1313,p1314,p1315,p1316,p1317,p1318,p1319,p1320,p1321,p1322,p1323,p1324,p1325,p1326,p1327,p1328,p1329,p1330,p1331,p1332,p1333,p1334,p1335,p1336,p1337,p1338,p1339,p1340,p1341,p1342,p1343,p1344,p1345,p1346,p1347,p1348,p1349,p1350,p1351,p1352,p1353,p1354,p1355,p1356,p1357,p1358,p1359,p1360,p1361,p1362,p1363,p1364,p1365,p1366,p1367,p1368,p1369,p1370,p1371,p1372,p1373,p1374,p1375,p1376,p1377,p1378,p1379,p1380,p1381,p1382,p1383,p1384,p1385,p1386,p1387,p1388,p1389,p1390,p1391,p1392,p1393,p1394,p1395,p1396,p1397,p1398,p1399,p1400,p1401,p1402,p1403,p1404,p1405,p1406,p1407,p1408,p1409,p1410,p1411,p1412,p1413,p1414,p1415,p1416,p1417,p1418,p1419,p1420,p1421,p1422,p1423,p1424,p1425,p1426,p1427,p1428,p1429,p1430,p1431,p1432,p1433,p1434,p1435,p1436,p1437,p1438,p1439,p1440,p1441,p1442,p1443,p1444,p1445,p1446,p1447,p1448,p1449,p1450,p1451,p1452,p1453,p1454,p1455,p1456,p1457,p1458,p1459,p1460,p1461,p1462,p1463,p1464,p1465,p1466,p1467,p1468,p1469,p1470,p1471,p1472,p1473,p1474,p1475,p1476,p1477,p1478,p1479,p1480,p1481,p1482,p1483,p1484,p1485,p1486,p1487,p1488,p1489,p1490,p1491,p1492,p1493,p1494,p1495,p1496,p1497,p1498,p1499,p1500,p1501,p1502,p1503,p1504,p1505,p1506,p1507,p1508,p1509,p1510,p1511,p1512,p1513,p1514,p1515,p1516,p1517,p1518,p1519,p1520,p1521,p1522,p1523,p1524,p1525,p1526,p1527,p1528,p1529,p1530,p1531,p1532,p1533,p1534,p1535,p1536,p1537,p1538,p1539,p1540,p1541,p1542,p1543,p1544,p1545,p1546,p1547,p1548,p1549,p1550,p1551,p1552,p1553,p1554,p1555,p1556,p1557,p1558,p1559,p1560,p1561,p1562,p1563,p1564,p1565,p1566,p1567,p1568,p1569,p1570,p1571,p1572,p1573,p1574,p1575,p1576,p1577,p1578,p1579,p1580,p1581,p1582,p1583,p1584,p1585,p1586,p1587,p1588,p1589,p1590,p1591,p1592,p1593,p1594,p1595,p1596,p1597,p1598,p1599,p1600,p1601,p1602,p1603,p1604,p1605,p1606,p1607,p1608,p1609,p1610,p1611,p1612,p1613,p1614,p1615,p1616,p1617,p1618,p1619,p1620,p1621,p1622,p1623,p1624,p1625,p1626,p1627,p1628,p1629,p1630,p1631,p1632,p1633,p1634,p1635,p1636,p1637,p1638,p1639,p1640,p1641,p1642,p1643,p1644,p1645,p1646,p1647,p1648,p1649,p1650,p1651,p1652,p1653,p1654,p1655,p1656,p1657,p1658,p1659,p1660,p1661,p1662,p1663,p1664,p1665,p1666,p1667,p1668,p1669,p1670,p1671,p1672,p1673,p1674,p1675,p1676,p1677,p1678,p1679,p1680,p1681,p1682,p1683,p1684,p1685,p1686,p1687,p1688,p1689,p1690,p1691,p1692,p1693,p1694,p1695,p1696,p1697,p1698,p1699,p1700,p1701,p1702,p1703,p1704,p1705,p1706,p1707,p1708,p1709,p1710,p1711,p1712,p1713,p1714,p1715,p1716,p1717,p1718,p1719,p1720,p1721,p1722,p1723,p1724,p1725,p1726,p1727,p1728,p1729,p1730,p1731,p1732,p1733,p1734,p1735,p1736,p1737,p1738,p1739,p1740,p1741,p1742,p1743,p1744,p1745,p1746,p1747,p1748,p1749,p1750,p1751,p1752,p1753,p1754,p1755,p1756,p1757,p1758,p1759,p1760,p1761,p1762,p1763,p1764,p1765,p1766,p1767,p1768,p1769,p1770,p1771,p1772,p1773,p1774,p1775,p1776,p1777,p1778,p1779,p1780,p1781,p1782,p1783,p1784,p1785,p1786,p1787,p1788,p1789,p1790,p1791,p1792,p1793,p1794,p1795,p1796,p1797,p1798,p1799,p1800,p1801,p1802,p1803,p1804,p1805,p1806,p1807,p1808,p1809,p1810,p1811,p1812,p1813,p1814,p1815,p1816,p1817,p1818,p1819,p1820,p1821,p1822,p1823,p1824,p1825,p1826,p1827,p1828,p1829,p1830,p1831,p1832,p1833,p1834,p1835,p1836,p1837,p1838,p1839,p1840,p1841,p1842,p1843,p1844,p1845,p1846,p1847,p1848,p1849,p1850,p1851,p1852,p1853,p1854,p1855,p1856,p1857,p1858,p1859,p1860,p1861,p1862,p1863,p1864,p1865,p1866,p1867,p1868,p1869,p1870,p1871,p1872,p1873,p1874,p1875,p1876,p1877,p1878,p1879,p1880,p1881,p1882,p1883,p1884,p1885,p1886,p1887,p1888,p1889,p1890,p1891,p1892,p1893,p1894,p1895,p1896,p1897,p1898,p1899,p1900,p1901,p1902,p1903,p1904,p1905,p1906,p1907,p1908,p1909,p1910,p1911,p1912,p1913,p1914,p1915,p1916,p1917,p1918,p1919,p1920,p1921,p1922,p1923,p1924,p1925,p1926,p1927,p1928,p1929,p1930,p1931,p1932,p1933,p1934,p1935,p1936,p1937,p1938,p1939,p1940,p1941,p1942,p1943,p1944,p1945,p1946,p1947,p1948,p1949,p1950,p1951,p1952,p1953,p1954,p1955,p1956,p1957,p1958,p1959,p1960,p1961,p1962,p1963,p1964,p1965,p1966,p1967,p1968,p1969,p1970,p1971,p1972,p1973,p1974,p1975,p1976,p1977,p1978,p1979,p1980,p1981,p1982,p1983,p1984,p1985,p1986,p1987,p1988,p1989,p1990,p1991,p1992,p1993,p1994,p1995,p1996,p1997,p1998,p1999,p2000,p2001,p2002,p2003,p2004,p2005,p2006,p2007,p2008,p2009,p2010,p2011,p2012,p2013,p2014,p2015,p2016,p2017,p2018,p2019,p2020,p2021,p2022,p2023,p2024,p2025,p2026,p2027,p2028,p2029,p2030,p2031,p2032,p2033,p2034,p2035,p2036,p2037,p2038,p2039,p2040,p2041,p2042,p2043,p2044,p2045,p2046,p2047,p2048,p2049,p2050,p2051,p2052,p2053,p2054,p2055,p2056,p2057,p2058,p2059,p2060,p2061,p2062,p2063,p2064,p2065,p2066,p2067,p2068,p2069,p2070,p2071,p2072,p2073,p2074,p2075,p2076,p2077,p2078,p2079,p2080,p2081,p2082,p2083,p2084,p2085,p2086,p2087,p2088,p2089,p2090,p2091,p2092,p2093,p2094,p2095,p2096,p2097,p2098,p2099,p2100,p2101,p2102,p2103,p2104,p2105,p2106,p2107,p2108,p2109,p2110,p2111,p2112,p2113,p2114,p2115,p2116,p2117,p2118,p2119,p2120,p2121,p2122,p2123,p2124,p2125,p2126,p2127,p2128,p2129,p2130,p2131,p2132,p2133,p2134,p2135,p2136,p2137,p2138,p2139,p2140,p2141,p2142,p2143,p2144,p2145,p2146,p2147,p2148,p2149,p2150,p2151,p2152,p2153,p2154,p2155,p2156,p2157,p2158,p2159,p2160,p2161,p2162,p2163,p2164,p2165,p2166,p2167,p2168,p2169,p2170,p2171,p2172,p2173,p2174,p2175,p2176,p2177,p2178,p2179,p2180,p2181,p2182,p2183,p2184,p2185,p2186,p2187,p2188,p2189,p2190,p2191,p2192,p2193,p2194,p2195,p2196,p2197,p2198,p2199,p2200,p2201,p2202,p2203,p2204,p2205,p2206,p2207,p2208,p2209,p2210,p2211,p2212,p2213,p2214,p2215,p2216,p2217,p2218,p2219,p2220,p2221,p2222,p2223,p2224,p2225,p2226,p2227,p2228,p2229,p2230,p2231,p2232,p2233,p2234,p2235,p2236,p2237,p2238,p2239,p2240,p2241,p2242,p2243,p2244,p2245,p2246,p2247,p2248,p2249,p2250,p2251,p2252,p2253,p2254,p2255,p2256,p2257,p2258,p2259,p2260,p2261,p2262,p2263,p2264,p2265,p2266,p2267,p2268,p2269,p2270,p2271,p2272,p2273,p2274,p2275,p2276,p2277,p2278,p2279,p2280,p2281,p2282,p2283,p2284,p2285,p2286,p2287,p2288,p2289,p2290,p2291,p2292,p2293,p2294,p2295,p2296,p2297,p2298,p2299,p2300,p2301,p2302,p2303,p2304,p2305,p2306,p2307,p2308,p2309,p2310,p2311,p2312,p2313,p2314,p2315,p2316,p2317,p2318,p2319,p2320,p2321,p2322,p2323,p2324,p2325,p2326,p2327,p2328,p2329,p2330,p2331,p2332,p2333,p2334,p2335,p2336,p2337,p2338,p2339,p2340,p2341,p2342,p2343,p2344,p2345,p2346,p2347,p2348,p2349,p2350,p2351,p2352,p2353,p2354,p2355,p2356,p2357,p2358,p2359,p2360,p2361,p2362,p2363,p2364,p2365,p2366,p2367,p2368,p2369,p2370,p2371,p2372,p2373,p2374,p2375,p2376,p2377,p2378,p2379,p2380,p2381,p2382,p2383,p2384,p2385,p2386,p2387,p2388,p2389,p2390,p2391,p2392,p2393,p2394,p2395,p2396,p2397,p2398,p2399,p2400,p2401,p2402,p2403,p2404,p2405,p2406,p2407,p2408,p2409,p2410,p2411,p2412,p2413,p2414,p2415,p2416,p2417,p2418,p2419,p2420,p2421,p2422,p2423,p2424,p2425,p2426,p2427,p2428,p2429,p2430,p2431,p2432,p2433,p2434,p2435,p2436,p2437,p2438,p2439,p2440,p2441,p2442,p2443,p2444,p2445,p2446,p2447,p2448,p2449,p2450,p2451,p2452,p2453,p2454,p2455,p2456,p2457,p2458,p2459,p2460,p2461,p2462,p2463,p2464,p2465,p2466,p2467,p2468,p2469,p2470,p2471,p2472,p2473,p2474,p2475,p2476,p2477,p2478,p2479,p2480,p2481,p2482,p2483,p2484,p2485,p2486,p2487,p2488,p2489,p2490,p2491,p2492,p2493,p2494,p2495,p2496,p2497,p2498,p2499,p2500,p2501,p2502,p2503,p2504,p2505,p2506,p2507,p2508,p2509,p2510,p2511,p2512,p2513,p2514,p2515,p2516,p2517,p2518,p2519,p2520,p2521,p2522,p2523,p2524,p2525,p2526,p2527,p2528,p2529,p2530,p2531,p2532,p2533,p2534,p2535,p2536,p2537,p2538,p2539,p2540,p2541,p2542,p2543,p2544,p2545,p2546,p2547,p2548,p2549,p2550,p2551,p2552,p2553,p2554,p2555,p2556,p2557,p2558,p2559,p2560,p2561,p2562,p2563,p2564,p2565,p2566,p2567,p2568,p2569,p2570,p2571,p2572,p2573,p2574,p2575,p2576,p2577,p2578,p2579,p2580,p2581,p2582,p2583,p2584,p2585,p2586,p2587,p2588,p2589,p2590,p2591,p2592,p2593,p2594,p2595,p2596,p2597,p2598,p2599,p2600,p2601,p2602,p2603,p2604,p2605,p2606,p2607,p2608,p2609,p2610,p2611,p2612,p2613,p2614,p2615,p2616,p2617,p2618,p2619,p2620,p2621,p2622,p2623,p2624,p2625,p2626,p2627,p2628,p2629,p2630,p2631,p2632,p2633,p2634,p2635,p2636,p2637,p2638,p2639,p2640,p2641,p2642,p2643,p2644,p2645,p2646,p2647,p2648,p2649,p2650,p2651,p2652,p2653,p2654,p2655,p2656,p2657,p2658,p2659,p2660,p2661,p2662,p2663,p2664,p2665,p2666,p2667,p2668,p2669,p2670,p2671,p2672,p2673,p2674,p2675,p2676,p2677,p2678,p2679,p2680,p2681,p2682,p2683,p2684,p2685,p2686,p2687,p2688,p2689,p2690,p2691,p2692,p2693,p2694,p2695,p2696,p2697,p2698,p2699,p2700,p2701,p2702,p2703,p2704,p2705,p2706,p2707,p2708,p2709,p2710,p2711,p2712,p2713,p2714,p2715,p2716,p2717,p2718,p2719,p2720,p2721,p2722,p2723,p2724,p2725,p2726,p2727,p2728,p2729,p2730,p2731,p2732,p2733,p2734,p2735,p2736,p2737,p2738,p2739,p2740,p2741,p2742,p2743,p2744,p2745,p2746,p2747,p2748,p2749,p2750,p2751,p2752,p2753,p2754,p2755,p2756,p2757,p2758,p2759,p2760,p2761,p2762,p2763,p2764,p2765,p2766,p2767,p2768,p2769,p2770,p2771,p2772,p2773,p2774,p2775,p2776,p2777,p2778,p2779,p2780,p2781,p2782,p2783,p2784,p2785,p2786,p2787,p2788,p2789,p2790,p2791,p2792,p2793,p2794,p2795,p2796,p2797,p2798,p2799,p2800,p2801,p2802,p2803,p2804,p2805,p2806,p2807,p2808,p2809,p2810,p2811,p2812,p2813,p2814,p2815,p2816,p2817,p2818,p2819,p2820,p2821,p2822,p2823,p2824,p2825,p2826,p2827,p2828,p2829,p2830,p2831,p2832,p2833,p2834,p2835,p2836,p2837,p2838,p2839,p2840,p2841,p2842,p2843,p2844,p2845,p2846,p2847,p2848,p2849,p2850,p2851,p2852,p2853,p2854,p2855,p2856,p2857,p2858,p2859,p2860,p2861,p2862,p2863,p2864,p2865,p2866,p2867,p2868,p2869,p2870,p2871,p2872,p2873,p2874,p2875,p2876,p2877,p2878,p2879,p2880,p2881,p2882,p2883,p2884,p2885,p2886,p2887,p2888,p2889,p2890,p2891,p2892,p2893,p2894,p2895,p2896,p2897,p2898,p2899,p2900,p2901,p2902,p2903,p2904,p2905,p2906,p2907,p2908,p2909,p2910,p2911,p2912,p2913,p2914,p2915,p2916,p2917,p2918,p2919,p2920,p2921,p2922,p2923,p2924,p2925,p2926,p2927,p2928,p2929,p2930,p2931,p2932,p2933,p2934,p2935,p2936,p2937,p2938,p2939,p2940,p2941,p2942,p2943,p2944,p2945,p2946,p2947,p2948,p2949,p2950,p2951,p2952,p2953,p2954,p2955,p2956,p2957,p2958,p2959,p2960,p2961,p2962,p2963,p2964,p2965,p2966,p2967,p2968,p2969,p2970,p2971,p2972,p2973,p2974,p2975,p2976,p2977,p2978,p2979,p2980,p2981,p2982,p2983,p2984,p2985,p2986,p2987,p2988,p2989,p2990,p2991,p2992,p2993,p2994,p2995,p2996,p2997,p2998,p2999,p3000,p3001,p3002,p3003,p3004,p3005,p3006,p3007,p3008,p3009,p3010,p3011,p3012,p3013,p3014,p3015,p3016,p3017,p3018,p3019,p3020,p3021,p3022,p3023,p3024,p3025,p3026,p3027,p3028,p3029,p3030,p3031,p3032,p3033,p3034,p3035,p3036,p3037,p3038,p3039,p3040,p3041,p3042,p3043,p3044,p3045,p3046,p3047,p3048,p3049,p3050,p3051,p3052,p3053,p3054,p3055,p3056,p3057,p3058,p3059,p3060,p3061,p3062,p3063,p3064,p3065,p3066,p3067,p3068,p3069,p3070,p3071,p3072,p3073,p3074,p3075,p3076,p3077,p3078,p3079,p3080,p3081,p3082,p3083,p3084,p3085,p3086,p3087,p3088,p3089,p3090,p3091,p3092,p3093,p3094,p3095,p3096,p3097,p3098,p3099,p3100,p3101,p3102,p3103,p3104,p3105,p3106,p3107,p3108,p3109,p3110,p3111,p3112,p3113,p3114,p3115,p3116,p3117,p3118,p3119,p3120,p3121,p3122,p3123;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_1_0,x[1],y[0]);
and and17(ip_1_1,x[1],y[1]);
and and18(ip_1_2,x[1],y[2]);
and and19(ip_1_3,x[1],y[3]);
and and20(ip_1_4,x[1],y[4]);
and and21(ip_1_5,x[1],y[5]);
and and22(ip_1_6,x[1],y[6]);
and and23(ip_1_7,x[1],y[7]);
and and24(ip_1_8,x[1],y[8]);
and and25(ip_1_9,x[1],y[9]);
and and26(ip_1_10,x[1],y[10]);
and and27(ip_1_11,x[1],y[11]);
and and28(ip_1_12,x[1],y[12]);
and and29(ip_1_13,x[1],y[13]);
and and30(ip_1_14,x[1],y[14]);
and and31(ip_1_15,x[1],y[15]);
and and32(ip_2_0,x[2],y[0]);
and and33(ip_2_1,x[2],y[1]);
and and34(ip_2_2,x[2],y[2]);
and and35(ip_2_3,x[2],y[3]);
and and36(ip_2_4,x[2],y[4]);
and and37(ip_2_5,x[2],y[5]);
and and38(ip_2_6,x[2],y[6]);
and and39(ip_2_7,x[2],y[7]);
and and40(ip_2_8,x[2],y[8]);
and and41(ip_2_9,x[2],y[9]);
and and42(ip_2_10,x[2],y[10]);
and and43(ip_2_11,x[2],y[11]);
and and44(ip_2_12,x[2],y[12]);
and and45(ip_2_13,x[2],y[13]);
and and46(ip_2_14,x[2],y[14]);
and and47(ip_2_15,x[2],y[15]);
and and48(ip_3_0,x[3],y[0]);
and and49(ip_3_1,x[3],y[1]);
and and50(ip_3_2,x[3],y[2]);
and and51(ip_3_3,x[3],y[3]);
and and52(ip_3_4,x[3],y[4]);
and and53(ip_3_5,x[3],y[5]);
and and54(ip_3_6,x[3],y[6]);
and and55(ip_3_7,x[3],y[7]);
and and56(ip_3_8,x[3],y[8]);
and and57(ip_3_9,x[3],y[9]);
and and58(ip_3_10,x[3],y[10]);
and and59(ip_3_11,x[3],y[11]);
and and60(ip_3_12,x[3],y[12]);
and and61(ip_3_13,x[3],y[13]);
and and62(ip_3_14,x[3],y[14]);
and and63(ip_3_15,x[3],y[15]);
and and64(ip_4_0,x[4],y[0]);
and and65(ip_4_1,x[4],y[1]);
and and66(ip_4_2,x[4],y[2]);
and and67(ip_4_3,x[4],y[3]);
and and68(ip_4_4,x[4],y[4]);
and and69(ip_4_5,x[4],y[5]);
and and70(ip_4_6,x[4],y[6]);
and and71(ip_4_7,x[4],y[7]);
and and72(ip_4_8,x[4],y[8]);
and and73(ip_4_9,x[4],y[9]);
and and74(ip_4_10,x[4],y[10]);
and and75(ip_4_11,x[4],y[11]);
and and76(ip_4_12,x[4],y[12]);
and and77(ip_4_13,x[4],y[13]);
and and78(ip_4_14,x[4],y[14]);
and and79(ip_4_15,x[4],y[15]);
and and80(ip_5_0,x[5],y[0]);
and and81(ip_5_1,x[5],y[1]);
and and82(ip_5_2,x[5],y[2]);
and and83(ip_5_3,x[5],y[3]);
and and84(ip_5_4,x[5],y[4]);
and and85(ip_5_5,x[5],y[5]);
and and86(ip_5_6,x[5],y[6]);
and and87(ip_5_7,x[5],y[7]);
and and88(ip_5_8,x[5],y[8]);
and and89(ip_5_9,x[5],y[9]);
and and90(ip_5_10,x[5],y[10]);
and and91(ip_5_11,x[5],y[11]);
and and92(ip_5_12,x[5],y[12]);
and and93(ip_5_13,x[5],y[13]);
and and94(ip_5_14,x[5],y[14]);
and and95(ip_5_15,x[5],y[15]);
and and96(ip_6_0,x[6],y[0]);
and and97(ip_6_1,x[6],y[1]);
and and98(ip_6_2,x[6],y[2]);
and and99(ip_6_3,x[6],y[3]);
and and100(ip_6_4,x[6],y[4]);
and and101(ip_6_5,x[6],y[5]);
and and102(ip_6_6,x[6],y[6]);
and and103(ip_6_7,x[6],y[7]);
and and104(ip_6_8,x[6],y[8]);
and and105(ip_6_9,x[6],y[9]);
and and106(ip_6_10,x[6],y[10]);
and and107(ip_6_11,x[6],y[11]);
and and108(ip_6_12,x[6],y[12]);
and and109(ip_6_13,x[6],y[13]);
and and110(ip_6_14,x[6],y[14]);
and and111(ip_6_15,x[6],y[15]);
and and112(ip_7_0,x[7],y[0]);
and and113(ip_7_1,x[7],y[1]);
and and114(ip_7_2,x[7],y[2]);
and and115(ip_7_3,x[7],y[3]);
and and116(ip_7_4,x[7],y[4]);
and and117(ip_7_5,x[7],y[5]);
and and118(ip_7_6,x[7],y[6]);
and and119(ip_7_7,x[7],y[7]);
and and120(ip_7_8,x[7],y[8]);
and and121(ip_7_9,x[7],y[9]);
and and122(ip_7_10,x[7],y[10]);
and and123(ip_7_11,x[7],y[11]);
and and124(ip_7_12,x[7],y[12]);
and and125(ip_7_13,x[7],y[13]);
and and126(ip_7_14,x[7],y[14]);
and and127(ip_7_15,x[7],y[15]);
and and128(ip_8_0,x[8],y[0]);
and and129(ip_8_1,x[8],y[1]);
and and130(ip_8_2,x[8],y[2]);
and and131(ip_8_3,x[8],y[3]);
and and132(ip_8_4,x[8],y[4]);
and and133(ip_8_5,x[8],y[5]);
and and134(ip_8_6,x[8],y[6]);
and and135(ip_8_7,x[8],y[7]);
and and136(ip_8_8,x[8],y[8]);
and and137(ip_8_9,x[8],y[9]);
and and138(ip_8_10,x[8],y[10]);
and and139(ip_8_11,x[8],y[11]);
and and140(ip_8_12,x[8],y[12]);
and and141(ip_8_13,x[8],y[13]);
and and142(ip_8_14,x[8],y[14]);
and and143(ip_8_15,x[8],y[15]);
and and144(ip_9_0,x[9],y[0]);
and and145(ip_9_1,x[9],y[1]);
and and146(ip_9_2,x[9],y[2]);
and and147(ip_9_3,x[9],y[3]);
and and148(ip_9_4,x[9],y[4]);
and and149(ip_9_5,x[9],y[5]);
and and150(ip_9_6,x[9],y[6]);
and and151(ip_9_7,x[9],y[7]);
and and152(ip_9_8,x[9],y[8]);
and and153(ip_9_9,x[9],y[9]);
and and154(ip_9_10,x[9],y[10]);
and and155(ip_9_11,x[9],y[11]);
and and156(ip_9_12,x[9],y[12]);
and and157(ip_9_13,x[9],y[13]);
and and158(ip_9_14,x[9],y[14]);
and and159(ip_9_15,x[9],y[15]);
and and160(ip_10_0,x[10],y[0]);
and and161(ip_10_1,x[10],y[1]);
and and162(ip_10_2,x[10],y[2]);
and and163(ip_10_3,x[10],y[3]);
and and164(ip_10_4,x[10],y[4]);
and and165(ip_10_5,x[10],y[5]);
and and166(ip_10_6,x[10],y[6]);
and and167(ip_10_7,x[10],y[7]);
and and168(ip_10_8,x[10],y[8]);
and and169(ip_10_9,x[10],y[9]);
and and170(ip_10_10,x[10],y[10]);
and and171(ip_10_11,x[10],y[11]);
and and172(ip_10_12,x[10],y[12]);
and and173(ip_10_13,x[10],y[13]);
and and174(ip_10_14,x[10],y[14]);
and and175(ip_10_15,x[10],y[15]);
and and176(ip_11_0,x[11],y[0]);
and and177(ip_11_1,x[11],y[1]);
and and178(ip_11_2,x[11],y[2]);
and and179(ip_11_3,x[11],y[3]);
and and180(ip_11_4,x[11],y[4]);
and and181(ip_11_5,x[11],y[5]);
and and182(ip_11_6,x[11],y[6]);
and and183(ip_11_7,x[11],y[7]);
and and184(ip_11_8,x[11],y[8]);
and and185(ip_11_9,x[11],y[9]);
and and186(ip_11_10,x[11],y[10]);
and and187(ip_11_11,x[11],y[11]);
and and188(ip_11_12,x[11],y[12]);
and and189(ip_11_13,x[11],y[13]);
and and190(ip_11_14,x[11],y[14]);
and and191(ip_11_15,x[11],y[15]);
and and192(ip_12_0,x[12],y[0]);
and and193(ip_12_1,x[12],y[1]);
and and194(ip_12_2,x[12],y[2]);
and and195(ip_12_3,x[12],y[3]);
and and196(ip_12_4,x[12],y[4]);
and and197(ip_12_5,x[12],y[5]);
and and198(ip_12_6,x[12],y[6]);
and and199(ip_12_7,x[12],y[7]);
and and200(ip_12_8,x[12],y[8]);
and and201(ip_12_9,x[12],y[9]);
and and202(ip_12_10,x[12],y[10]);
and and203(ip_12_11,x[12],y[11]);
and and204(ip_12_12,x[12],y[12]);
and and205(ip_12_13,x[12],y[13]);
and and206(ip_12_14,x[12],y[14]);
and and207(ip_12_15,x[12],y[15]);
and and208(ip_13_0,x[13],y[0]);
and and209(ip_13_1,x[13],y[1]);
and and210(ip_13_2,x[13],y[2]);
and and211(ip_13_3,x[13],y[3]);
and and212(ip_13_4,x[13],y[4]);
and and213(ip_13_5,x[13],y[5]);
and and214(ip_13_6,x[13],y[6]);
and and215(ip_13_7,x[13],y[7]);
and and216(ip_13_8,x[13],y[8]);
and and217(ip_13_9,x[13],y[9]);
and and218(ip_13_10,x[13],y[10]);
and and219(ip_13_11,x[13],y[11]);
and and220(ip_13_12,x[13],y[12]);
and and221(ip_13_13,x[13],y[13]);
and and222(ip_13_14,x[13],y[14]);
and and223(ip_13_15,x[13],y[15]);
and and224(ip_14_0,x[14],y[0]);
and and225(ip_14_1,x[14],y[1]);
and and226(ip_14_2,x[14],y[2]);
and and227(ip_14_3,x[14],y[3]);
and and228(ip_14_4,x[14],y[4]);
and and229(ip_14_5,x[14],y[5]);
and and230(ip_14_6,x[14],y[6]);
and and231(ip_14_7,x[14],y[7]);
and and232(ip_14_8,x[14],y[8]);
and and233(ip_14_9,x[14],y[9]);
and and234(ip_14_10,x[14],y[10]);
and and235(ip_14_11,x[14],y[11]);
and and236(ip_14_12,x[14],y[12]);
and and237(ip_14_13,x[14],y[13]);
and and238(ip_14_14,x[14],y[14]);
and and239(ip_14_15,x[14],y[15]);
and and240(ip_15_0,x[15],y[0]);
and and241(ip_15_1,x[15],y[1]);
and and242(ip_15_2,x[15],y[2]);
and and243(ip_15_3,x[15],y[3]);
and and244(ip_15_4,x[15],y[4]);
and and245(ip_15_5,x[15],y[5]);
and and246(ip_15_6,x[15],y[6]);
and and247(ip_15_7,x[15],y[7]);
and and248(ip_15_8,x[15],y[8]);
and and249(ip_15_9,x[15],y[9]);
and and250(ip_15_10,x[15],y[10]);
and and251(ip_15_11,x[15],y[11]);
and and252(ip_15_12,x[15],y[12]);
and and253(ip_15_13,x[15],y[13]);
and and254(ip_15_14,x[15],y[14]);
and and255(ip_15_15,x[15],y[15]);
HA ha0(ip_0_2,ip_1_1,p0,p1);
HA ha1(ip_0_3,ip_1_2,p2,p3);
HA ha2(ip_2_1,ip_3_0,p4,p5);
HA ha3(p0,p3,p6,p7);
HA ha4(ip_0_4,ip_1_3,p8,p9);
HA ha5(ip_2_2,ip_3_1,p10,p11);
HA ha6(ip_4_0,p11,p12,p13);
HA ha7(p2,p4,p14,p15);
HA ha8(p9,p13,p16,p17);
HA ha9(p15,p6,p18,p19);
HA ha10(ip_0_5,ip_1_4,p20,p21);
HA ha11(ip_2_3,ip_3_2,p22,p23);
HA ha12(ip_4_1,ip_5_0,p24,p25);
HA ha13(p10,p21,p26,p27);
HA ha14(p23,p25,p28,p29);
HA ha15(p8,p12,p30,p31);
HA ha16(p14,p27,p32,p33);
HA ha17(p29,p16,p34,p35);
HA ha18(p18,p31,p36,p37);
HA ha19(p33,p35,p38,p39);
HA ha20(ip_0_6,ip_1_5,p40,p41);
HA ha21(ip_2_4,ip_3_3,p42,p43);
HA ha22(ip_4_2,ip_5_1,p44,p45);
HA ha23(ip_6_0,p20,p46,p47);
HA ha24(p22,p24,p48,p49);
HA ha25(p41,p43,p50,p51);
HA ha26(p45,p26,p52,p53);
HA ha27(p28,p47,p54,p55);
HA ha28(p49,p51,p56,p57);
HA ha29(p30,p32,p58,p59);
HA ha30(p53,p55,p60,p61);
HA ha31(p57,p34,p62,p63);
HA ha32(p36,p59,p64,p65);
HA ha33(p61,p38,p66,p67);
HA ha34(p63,p65,p68,p69);
FA fa0(ip_0_7,ip_1_6,ip_2_5,p70,p71);
HA ha35(ip_3_4,ip_4_3,p72,p73);
HA ha36(ip_5_2,ip_6_1,p74,p75);
HA ha37(ip_7_0,p40,p76,p77);
HA ha38(p42,p44,p78,p79);
HA ha39(p73,p75,p80,p81);
HA ha40(p46,p48,p82,p83);
HA ha41(p50,p71,p84,p85);
HA ha42(p77,p79,p86,p87);
HA ha43(p81,p52,p88,p89);
HA ha44(p54,p56,p90,p91);
HA ha45(p83,p85,p92,p93);
HA ha46(p87,p58,p94,p95);
HA ha47(p60,p89,p96,p97);
HA ha48(p91,p93,p98,p99);
HA ha49(p62,p64,p100,p101);
HA ha50(p95,p97,p102,p103);
FA fa1(p99,p101,p103,p104,p105);
HA ha51(p66,p68,p106,p107);
HA ha52(ip_0_8,ip_1_7,p108,p109);
HA ha53(ip_2_6,ip_3_5,p110,p111);
HA ha54(ip_4_4,ip_5_3,p112,p113);
HA ha55(ip_6_2,ip_7_1,p114,p115);
HA ha56(ip_8_0,p109,p116,p117);
HA ha57(p111,p113,p118,p119);
HA ha58(p115,p72,p120,p121);
HA ha59(p74,p117,p122,p123);
HA ha60(p119,p121,p124,p125);
HA ha61(p76,p78,p126,p127);
HA ha62(p80,p123,p128,p129);
HA ha63(p125,p127,p130,p131);
HA ha64(p70,p82,p132,p133);
HA ha65(p84,p86,p134,p135);
HA ha66(p129,p131,p136,p137);
HA ha67(p133,p135,p138,p139);
HA ha68(p88,p90,p140,p141);
FA fa2(p92,p137,p139,p142,p143);
HA ha69(p141,p94,p144,p145);
HA ha70(p96,p98,p146,p147);
FA fa3(p100,p102,p145,p148,p149);
HA ha71(p147,p106,p150,p151);
HA ha72(p143,p149,p152,p153);
HA ha73(p151,p104,p154,p155);
HA ha74(ip_0_9,ip_1_8,p156,p157);
HA ha75(ip_2_7,ip_3_6,p158,p159);
HA ha76(ip_4_5,ip_5_4,p160,p161);
HA ha77(ip_6_3,ip_7_2,p162,p163);
HA ha78(ip_8_1,ip_9_0,p164,p165);
HA ha79(p108,p110,p166,p167);
FA fa4(p112,p114,p157,p168,p169);
HA ha80(p159,p161,p170,p171);
HA ha81(p163,p165,p172,p173);
HA ha82(p116,p118,p174,p175);
HA ha83(p120,p167,p176,p177);
HA ha84(p171,p173,p178,p179);
HA ha85(p122,p124,p180,p181);
HA ha86(p126,p169,p182,p183);
HA ha87(p175,p177,p184,p185);
FA fa5(p179,p128,p130,p186,p187);
HA ha88(p132,p134,p188,p189);
HA ha89(p181,p183,p190,p191);
FA fa6(p185,p136,p138,p192,p193);
HA ha90(p140,p189,p194,p195);
HA ha91(p191,p144,p196,p197);
HA ha92(p146,p187,p198,p199);
HA ha93(p195,p193,p200,p201);
HA ha94(p197,p199,p202,p203);
HA ha95(p142,p150,p204,p205);
HA ha96(p201,p203,p206,p207);
HA ha97(p148,p152,p208,p209);
HA ha98(p205,p207,p210,p211);
FA fa7(p154,p209,p211,p212,p213);
HA ha99(ip_0_10,ip_1_9,p214,p215);
HA ha100(ip_2_8,ip_3_7,p216,p217);
HA ha101(ip_4_6,ip_5_5,p218,p219);
HA ha102(ip_6_4,ip_7_3,p220,p221);
HA ha103(ip_8_2,ip_9_1,p222,p223);
HA ha104(ip_10_0,p156,p224,p225);
HA ha105(p158,p160,p226,p227);
HA ha106(p162,p164,p228,p229);
HA ha107(p215,p217,p230,p231);
FA fa8(p219,p221,p223,p232,p233);
HA ha108(p166,p170,p234,p235);
HA ha109(p172,p225,p236,p237);
HA ha110(p227,p229,p238,p239);
HA ha111(p231,p174,p240,p241);
FA fa9(p176,p178,p233,p242,p243);
HA ha112(p235,p237,p244,p245);
HA ha113(p239,p168,p246,p247);
HA ha114(p180,p182,p248,p249);
HA ha115(p184,p241,p250,p251);
HA ha116(p245,p188,p252,p253);
HA ha117(p190,p243,p254,p255);
HA ha118(p247,p249,p256,p257);
HA ha119(p251,p194,p258,p259);
HA ha120(p253,p255,p260,p261);
HA ha121(p257,p186,p262,p263);
HA ha122(p196,p198,p264,p265);
HA ha123(p259,p261,p266,p267);
HA ha124(p192,p200,p268,p269);
HA ha125(p202,p263,p270,p271);
HA ha126(p265,p267,p272,p273);
HA ha127(p204,p206,p274,p275);
FA fa10(p269,p271,p273,p276,p277);
HA ha128(p208,p210,p278,p279);
HA ha129(p275,p277,p280,p281);
HA ha130(p279,p281,p282,p283);
HA ha131(ip_0_11,ip_1_10,p284,p285);
HA ha132(ip_2_9,ip_3_8,p286,p287);
HA ha133(ip_4_7,ip_5_6,p288,p289);
HA ha134(ip_6_5,ip_7_4,p290,p291);
HA ha135(ip_8_3,ip_9_2,p292,p293);
HA ha136(ip_10_1,ip_11_0,p294,p295);
HA ha137(p214,p216,p296,p297);
HA ha138(p218,p220,p298,p299);
HA ha139(p222,p285,p300,p301);
HA ha140(p287,p289,p302,p303);
HA ha141(p291,p293,p304,p305);
HA ha142(p295,p224,p306,p307);
HA ha143(p226,p228,p308,p309);
HA ha144(p230,p297,p310,p311);
HA ha145(p299,p301,p312,p313);
FA fa11(p303,p305,p234,p314,p315);
HA ha146(p236,p238,p316,p317);
HA ha147(p307,p309,p318,p319);
HA ha148(p311,p313,p320,p321);
HA ha149(p232,p240,p322,p323);
HA ha150(p244,p315,p324,p325);
HA ha151(p317,p319,p326,p327);
HA ha152(p321,p246,p328,p329);
HA ha153(p248,p250,p330,p331);
HA ha154(p323,p325,p332,p333);
HA ha155(p327,p242,p334,p335);
HA ha156(p252,p254,p336,p337);
HA ha157(p256,p329,p338,p339);
HA ha158(p331,p333,p340,p341);
HA ha159(p258,p260,p342,p343);
HA ha160(p335,p337,p344,p345);
HA ha161(p339,p341,p346,p347);
HA ha162(p262,p264,p348,p349);
HA ha163(p266,p343,p350,p351);
HA ha164(p345,p347,p352,p353);
HA ha165(p268,p270,p354,p355);
HA ha166(p272,p349,p356,p357);
HA ha167(p351,p353,p358,p359);
FA fa12(p274,p355,p357,p360,p361);
HA ha168(p359,p278,p362,p363);
HA ha169(p276,p280,p364,p365);
HA ha170(p361,p363,p366,p367);
HA ha171(p282,p365,p368,p369);
HA ha172(ip_0_12,ip_1_11,p370,p371);
HA ha173(ip_2_10,ip_3_9,p372,p373);
HA ha174(ip_4_8,ip_5_7,p374,p375);
HA ha175(ip_6_6,ip_7_5,p376,p377);
HA ha176(ip_8_4,ip_9_3,p378,p379);
HA ha177(ip_10_2,ip_11_1,p380,p381);
FA fa13(ip_12_0,p284,p286,p382,p383);
HA ha178(p288,p290,p384,p385);
HA ha179(p292,p294,p386,p387);
HA ha180(p371,p373,p388,p389);
HA ha181(p375,p377,p390,p391);
HA ha182(p379,p381,p392,p393);
HA ha183(p296,p298,p394,p395);
HA ha184(p300,p302,p396,p397);
HA ha185(p304,p385,p398,p399);
FA fa14(p387,p389,p391,p400,p401);
HA ha186(p393,p306,p402,p403);
HA ha187(p308,p310,p404,p405);
HA ha188(p312,p383,p406,p407);
HA ha189(p395,p397,p408,p409);
HA ha190(p399,p316,p410,p411);
HA ha191(p318,p320,p412,p413);
HA ha192(p401,p403,p414,p415);
HA ha193(p405,p407,p416,p417);
HA ha194(p409,p314,p418,p419);
FA fa15(p322,p324,p326,p420,p421);
HA ha195(p411,p413,p422,p423);
HA ha196(p415,p417,p424,p425);
HA ha197(p328,p330,p426,p427);
FA fa16(p332,p419,p423,p428,p429);
HA ha198(p425,p334,p430,p431);
HA ha199(p336,p338,p432,p433);
HA ha200(p340,p421,p434,p435);
HA ha201(p427,p342,p436,p437);
HA ha202(p344,p346,p438,p439);
HA ha203(p429,p431,p440,p441);
HA ha204(p433,p435,p442,p443);
FA fa17(p348,p350,p352,p444,p445);
HA ha205(p437,p439,p446,p447);
HA ha206(p441,p443,p448,p449);
FA fa18(p354,p356,p358,p450,p451);
HA ha207(p447,p449,p452,p453);
HA ha208(p445,p453,p454,p455);
HA ha209(p362,p451,p456,p457);
HA ha210(p455,p360,p458,p459);
HA ha211(p364,p366,p460,p461);
HA ha212(p457,p368,p462,p463);
HA ha213(p459,p461,p464,p465);
FA fa19(ip_0_13,ip_1_12,ip_2_11,p466,p467);
HA ha214(ip_3_10,ip_4_9,p468,p469);
HA ha215(ip_5_8,ip_6_7,p470,p471);
HA ha216(ip_7_6,ip_8_5,p472,p473);
HA ha217(ip_9_4,ip_10_3,p474,p475);
HA ha218(ip_11_2,ip_12_1,p476,p477);
HA ha219(ip_13_0,p370,p478,p479);
HA ha220(p372,p374,p480,p481);
HA ha221(p376,p378,p482,p483);
HA ha222(p380,p469,p484,p485);
HA ha223(p471,p473,p486,p487);
HA ha224(p475,p477,p488,p489);
HA ha225(p384,p386,p490,p491);
HA ha226(p388,p390,p492,p493);
HA ha227(p392,p467,p494,p495);
HA ha228(p479,p481,p496,p497);
FA fa20(p483,p485,p487,p498,p499);
HA ha229(p489,p394,p500,p501);
HA ha230(p396,p398,p502,p503);
HA ha231(p491,p493,p504,p505);
HA ha232(p495,p497,p506,p507);
HA ha233(p382,p402,p508,p509);
HA ha234(p404,p406,p510,p511);
HA ha235(p408,p499,p512,p513);
HA ha236(p501,p503,p514,p515);
HA ha237(p505,p507,p516,p517);
HA ha238(p400,p410,p518,p519);
HA ha239(p412,p414,p520,p521);
HA ha240(p416,p509,p522,p523);
HA ha241(p511,p513,p524,p525);
HA ha242(p515,p517,p526,p527);
HA ha243(p418,p422,p528,p529);
HA ha244(p424,p519,p530,p531);
HA ha245(p521,p523,p532,p533);
HA ha246(p525,p527,p534,p535);
HA ha247(p426,p529,p536,p537);
HA ha248(p531,p533,p538,p539);
HA ha249(p535,p420,p540,p541);
HA ha250(p430,p432,p542,p543);
HA ha251(p434,p537,p544,p545);
HA ha252(p539,p428,p546,p547);
HA ha253(p436,p438,p548,p549);
HA ha254(p440,p442,p550,p551);
HA ha255(p541,p543,p552,p553);
HA ha256(p545,p446,p554,p555);
HA ha257(p448,p547,p556,p557);
FA fa21(p549,p551,p553,p558,p559);
FA fa22(p452,p555,p557,p560,p561);
HA ha258(p444,p454,p562,p563);
HA ha259(p559,p450,p564,p565);
HA ha260(p456,p561,p566,p567);
HA ha261(p563,p458,p568,p569);
HA ha262(p460,p565,p570,p571);
HA ha263(p567,p462,p572,p573);
HA ha264(p464,p569,p574,p575);
FA fa23(p571,p573,p575,p576,p577);
HA ha265(ip_0_14,ip_1_13,p578,p579);
HA ha266(ip_2_12,ip_3_11,p580,p581);
HA ha267(ip_4_10,ip_5_9,p582,p583);
HA ha268(ip_6_8,ip_7_7,p584,p585);
HA ha269(ip_8_6,ip_9_5,p586,p587);
HA ha270(ip_10_4,ip_11_3,p588,p589);
FA fa24(ip_12_2,ip_13_1,ip_14_0,p590,p591);
HA ha271(p468,p470,p592,p593);
HA ha272(p472,p474,p594,p595);
HA ha273(p476,p579,p596,p597);
HA ha274(p581,p583,p598,p599);
HA ha275(p585,p587,p600,p601);
HA ha276(p589,p478,p602,p603);
HA ha277(p480,p482,p604,p605);
HA ha278(p484,p486,p606,p607);
HA ha279(p488,p591,p608,p609);
FA fa25(p593,p595,p597,p610,p611);
HA ha280(p599,p601,p612,p613);
FA fa26(p466,p490,p492,p614,p615);
HA ha281(p494,p496,p616,p617);
FA fa27(p603,p605,p607,p618,p619);
HA ha282(p609,p613,p620,p621);
HA ha283(p500,p502,p622,p623);
HA ha284(p504,p506,p624,p625);
HA ha285(p611,p617,p626,p627);
HA ha286(p621,p498,p628,p629);
HA ha287(p508,p510,p630,p631);
HA ha288(p512,p514,p632,p633);
HA ha289(p516,p615,p634,p635);
HA ha290(p619,p623,p636,p637);
HA ha291(p625,p627,p638,p639);
HA ha292(p518,p520,p640,p641);
HA ha293(p522,p524,p642,p643);
HA ha294(p526,p629,p644,p645);
HA ha295(p631,p633,p646,p647);
HA ha296(p635,p637,p648,p649);
HA ha297(p639,p528,p650,p651);
HA ha298(p530,p532,p652,p653);
HA ha299(p534,p641,p654,p655);
HA ha300(p643,p645,p656,p657);
HA ha301(p647,p649,p658,p659);
HA ha302(p536,p538,p660,p661);
HA ha303(p651,p653,p662,p663);
HA ha304(p655,p657,p664,p665);
HA ha305(p659,p540,p666,p667);
HA ha306(p542,p544,p668,p669);
HA ha307(p661,p663,p670,p671);
HA ha308(p665,p546,p672,p673);
HA ha309(p548,p550,p674,p675);
HA ha310(p552,p667,p676,p677);
HA ha311(p669,p671,p678,p679);
HA ha312(p554,p556,p680,p681);
HA ha313(p673,p675,p682,p683);
HA ha314(p677,p679,p684,p685);
HA ha315(p681,p683,p686,p687);
HA ha316(p685,p558,p688,p689);
HA ha317(p562,p687,p690,p691);
HA ha318(p560,p564,p692,p693);
HA ha319(p566,p689,p694,p695);
HA ha320(p691,p568,p696,p697);
HA ha321(p570,p693,p698,p699);
HA ha322(p695,p572,p700,p701);
HA ha323(p574,p697,p702,p703);
HA ha324(p699,p701,p704,p705);
HA ha325(p703,p705,p706,p707);
HA ha326(ip_0_15,ip_1_14,p708,p709);
HA ha327(ip_2_13,ip_3_12,p710,p711);
HA ha328(ip_4_11,ip_5_10,p712,p713);
FA fa28(ip_6_9,ip_7_8,ip_8_7,p714,p715);
HA ha329(ip_9_6,ip_10_5,p716,p717);
HA ha330(ip_11_4,ip_12_3,p718,p719);
HA ha331(ip_13_2,ip_14_1,p720,p721);
HA ha332(ip_15_0,p578,p722,p723);
HA ha333(p580,p582,p724,p725);
HA ha334(p584,p586,p726,p727);
HA ha335(p588,p709,p728,p729);
HA ha336(p711,p713,p730,p731);
HA ha337(p717,p719,p732,p733);
HA ha338(p721,p592,p734,p735);
HA ha339(p594,p596,p736,p737);
FA fa29(p598,p600,p715,p738,p739);
HA ha340(p723,p725,p740,p741);
HA ha341(p727,p729,p742,p743);
FA fa30(p731,p733,p590,p744,p745);
HA ha342(p602,p604,p746,p747);
HA ha343(p606,p608,p748,p749);
HA ha344(p612,p735,p750,p751);
HA ha345(p737,p741,p752,p753);
HA ha346(p743,p616,p754,p755);
HA ha347(p620,p739,p756,p757);
HA ha348(p745,p747,p758,p759);
HA ha349(p749,p751,p760,p761);
HA ha350(p753,p610,p762,p763);
HA ha351(p622,p624,p764,p765);
HA ha352(p626,p755,p766,p767);
HA ha353(p757,p759,p768,p769);
HA ha354(p761,p614,p770,p771);
HA ha355(p618,p628,p772,p773);
HA ha356(p630,p632,p774,p775);
HA ha357(p634,p636,p776,p777);
HA ha358(p638,p763,p778,p779);
HA ha359(p765,p767,p780,p781);
HA ha360(p769,p640,p782,p783);
HA ha361(p642,p644,p784,p785);
HA ha362(p646,p648,p786,p787);
HA ha363(p771,p773,p788,p789);
HA ha364(p775,p777,p790,p791);
HA ha365(p779,p781,p792,p793);
HA ha366(p650,p652,p794,p795);
HA ha367(p654,p656,p796,p797);
HA ha368(p658,p783,p798,p799);
HA ha369(p785,p787,p800,p801);
HA ha370(p789,p791,p802,p803);
HA ha371(p793,p660,p804,p805);
HA ha372(p662,p664,p806,p807);
HA ha373(p795,p797,p808,p809);
HA ha374(p799,p801,p810,p811);
HA ha375(p803,p666,p812,p813);
HA ha376(p668,p670,p814,p815);
FA fa31(p805,p807,p809,p816,p817);
HA ha377(p811,p672,p818,p819);
HA ha378(p674,p676,p820,p821);
HA ha379(p678,p813,p822,p823);
HA ha380(p815,p680,p824,p825);
HA ha381(p682,p684,p826,p827);
HA ha382(p817,p819,p828,p829);
HA ha383(p821,p823,p830,p831);
HA ha384(p686,p825,p832,p833);
HA ha385(p827,p829,p834,p835);
HA ha386(p831,p688,p836,p837);
FA fa32(p690,p833,p835,p838,p839);
HA ha387(p692,p694,p840,p841);
HA ha388(p837,p696,p842,p843);
HA ha389(p698,p839,p844,p845);
HA ha390(p841,p700,p846,p847);
HA ha391(p702,p843,p848,p849);
HA ha392(p845,p704,p850,p851);
HA ha393(p847,p849,p852,p853);
FA fa33(p706,p851,p853,p854,p855);
HA ha394(ip_1_15,ip_2_14,p856,p857);
HA ha395(ip_3_13,ip_4_12,p858,p859);
HA ha396(ip_5_11,ip_6_10,p860,p861);
HA ha397(ip_7_9,ip_8_8,p862,p863);
HA ha398(ip_9_7,ip_10_6,p864,p865);
HA ha399(ip_11_5,ip_12_4,p866,p867);
HA ha400(ip_13_3,ip_14_2,p868,p869);
HA ha401(ip_15_1,p708,p870,p871);
HA ha402(p710,p712,p872,p873);
HA ha403(p716,p718,p874,p875);
HA ha404(p720,p857,p876,p877);
HA ha405(p859,p861,p878,p879);
HA ha406(p863,p865,p880,p881);
HA ha407(p867,p869,p882,p883);
HA ha408(p722,p724,p884,p885);
FA fa34(p726,p728,p730,p886,p887);
HA ha409(p732,p871,p888,p889);
HA ha410(p873,p875,p890,p891);
HA ha411(p877,p879,p892,p893);
HA ha412(p881,p883,p894,p895);
FA fa35(p714,p734,p736,p896,p897);
HA ha413(p740,p742,p898,p899);
HA ha414(p885,p889,p900,p901);
HA ha415(p891,p893,p902,p903);
HA ha416(p895,p746,p904,p905);
HA ha417(p748,p750,p906,p907);
HA ha418(p752,p887,p908,p909);
HA ha419(p899,p901,p910,p911);
HA ha420(p903,p738,p912,p913);
HA ha421(p744,p754,p914,p915);
HA ha422(p756,p758,p916,p917);
HA ha423(p760,p897,p918,p919);
HA ha424(p905,p907,p920,p921);
HA ha425(p909,p911,p922,p923);
HA ha426(p762,p764,p924,p925);
HA ha427(p766,p768,p926,p927);
HA ha428(p913,p915,p928,p929);
HA ha429(p917,p919,p930,p931);
HA ha430(p921,p923,p932,p933);
HA ha431(p770,p772,p934,p935);
HA ha432(p774,p776,p936,p937);
HA ha433(p778,p780,p938,p939);
HA ha434(p925,p927,p940,p941);
HA ha435(p929,p931,p942,p943);
HA ha436(p933,p782,p944,p945);
HA ha437(p784,p786,p946,p947);
HA ha438(p788,p790,p948,p949);
HA ha439(p792,p935,p950,p951);
HA ha440(p937,p939,p952,p953);
HA ha441(p941,p943,p954,p955);
HA ha442(p794,p796,p956,p957);
HA ha443(p798,p800,p958,p959);
HA ha444(p802,p945,p960,p961);
HA ha445(p947,p949,p962,p963);
HA ha446(p951,p953,p964,p965);
HA ha447(p955,p804,p966,p967);
HA ha448(p806,p808,p968,p969);
HA ha449(p810,p957,p970,p971);
HA ha450(p959,p961,p972,p973);
HA ha451(p963,p965,p974,p975);
HA ha452(p812,p814,p976,p977);
HA ha453(p967,p969,p978,p979);
HA ha454(p971,p973,p980,p981);
HA ha455(p975,p818,p982,p983);
HA ha456(p820,p822,p984,p985);
HA ha457(p977,p979,p986,p987);
HA ha458(p981,p816,p988,p989);
HA ha459(p824,p826,p990,p991);
HA ha460(p828,p830,p992,p993);
HA ha461(p983,p985,p994,p995);
HA ha462(p987,p832,p996,p997);
HA ha463(p834,p989,p998,p999);
HA ha464(p991,p993,p1000,p1001);
HA ha465(p995,p1001,p1002,p1003);
HA ha466(p836,p997,p1004,p1005);
HA ha467(p999,p1003,p1006,p1007);
HA ha468(p1005,p840,p1008,p1009);
HA ha469(p1007,p1009,p1010,p1011);
HA ha470(p838,p842,p1012,p1013);
HA ha471(p844,p1011,p1014,p1015);
HA ha472(p1013,p846,p1016,p1017);
HA ha473(p848,p1015,p1018,p1019);
HA ha474(p1017,p850,p1020,p1021);
HA ha475(p852,p1019,p1022,p1023);
HA ha476(p1021,p1023,p1024,p1025);
FA fa36(ip_2_15,ip_3_14,ip_4_13,p1026,p1027);
HA ha477(ip_5_12,ip_6_11,p1028,p1029);
HA ha478(ip_7_10,ip_8_9,p1030,p1031);
HA ha479(ip_9_8,ip_10_7,p1032,p1033);
HA ha480(ip_11_6,ip_12_5,p1034,p1035);
HA ha481(ip_13_4,ip_14_3,p1036,p1037);
HA ha482(ip_15_2,p1029,p1038,p1039);
FA fa37(p1031,p1033,p1035,p1040,p1041);
HA ha483(p1037,p856,p1042,p1043);
HA ha484(p858,p860,p1044,p1045);
HA ha485(p862,p864,p1046,p1047);
HA ha486(p866,p868,p1048,p1049);
HA ha487(p1027,p1039,p1050,p1051);
HA ha488(p1043,p1045,p1052,p1053);
HA ha489(p1047,p1049,p1054,p1055);
HA ha490(p870,p872,p1056,p1057);
HA ha491(p874,p876,p1058,p1059);
HA ha492(p878,p880,p1060,p1061);
HA ha493(p882,p1041,p1062,p1063);
HA ha494(p1051,p1053,p1064,p1065);
HA ha495(p1055,p1057,p1066,p1067);
HA ha496(p1059,p1061,p1068,p1069);
HA ha497(p884,p888,p1070,p1071);
HA ha498(p890,p892,p1072,p1073);
HA ha499(p894,p1063,p1074,p1075);
HA ha500(p1065,p1067,p1076,p1077);
HA ha501(p1069,p1071,p1078,p1079);
HA ha502(p1073,p898,p1080,p1081);
HA ha503(p900,p902,p1082,p1083);
HA ha504(p1075,p1077,p1084,p1085);
HA ha505(p1079,p1081,p1086,p1087);
HA ha506(p1083,p886,p1088,p1089);
HA ha507(p904,p906,p1090,p1091);
FA fa38(p908,p910,p1085,p1092,p1093);
HA ha508(p1087,p1089,p1094,p1095);
HA ha509(p1091,p896,p1096,p1097);
HA ha510(p912,p914,p1098,p1099);
HA ha511(p916,p918,p1100,p1101);
HA ha512(p920,p922,p1102,p1103);
HA ha513(p1093,p1095,p1104,p1105);
FA fa39(p1097,p1099,p1101,p1106,p1107);
FA fa40(p1103,p924,p926,p1108,p1109);
HA ha514(p928,p930,p1110,p1111);
HA ha515(p932,p1105,p1112,p1113);
HA ha516(p1111,p934,p1114,p1115);
HA ha517(p936,p938,p1116,p1117);
HA ha518(p940,p942,p1118,p1119);
HA ha519(p1107,p1109,p1120,p1121);
HA ha520(p1113,p1115,p1122,p1123);
HA ha521(p1117,p1119,p1124,p1125);
HA ha522(p944,p946,p1126,p1127);
HA ha523(p948,p950,p1128,p1129);
HA ha524(p952,p954,p1130,p1131);
HA ha525(p1121,p1123,p1132,p1133);
HA ha526(p1125,p1127,p1134,p1135);
HA ha527(p1129,p1131,p1136,p1137);
HA ha528(p956,p958,p1138,p1139);
HA ha529(p960,p962,p1140,p1141);
HA ha530(p964,p1133,p1142,p1143);
HA ha531(p1135,p1137,p1144,p1145);
HA ha532(p1139,p1141,p1146,p1147);
HA ha533(p966,p968,p1148,p1149);
HA ha534(p970,p972,p1150,p1151);
HA ha535(p974,p1143,p1152,p1153);
HA ha536(p1145,p1147,p1154,p1155);
HA ha537(p1149,p1151,p1156,p1157);
HA ha538(p976,p978,p1158,p1159);
HA ha539(p980,p1153,p1160,p1161);
HA ha540(p1155,p1157,p1162,p1163);
HA ha541(p1159,p982,p1164,p1165);
HA ha542(p984,p986,p1166,p1167);
HA ha543(p1161,p1163,p1168,p1169);
HA ha544(p1165,p1167,p1170,p1171);
HA ha545(p988,p990,p1172,p1173);
HA ha546(p992,p994,p1174,p1175);
HA ha547(p1000,p1169,p1176,p1177);
HA ha548(p1171,p1173,p1178,p1179);
HA ha549(p1175,p996,p1180,p1181);
HA ha550(p998,p1002,p1182,p1183);
HA ha551(p1004,p1177,p1184,p1185);
HA ha552(p1179,p1181,p1186,p1187);
FA fa41(p1006,p1008,p1183,p1188,p1189);
HA ha553(p1185,p1187,p1190,p1191);
HA ha554(p1010,p1012,p1192,p1193);
HA ha555(p1191,p1014,p1194,p1195);
HA ha556(p1016,p1189,p1196,p1197);
HA ha557(p1193,p1018,p1198,p1199);
HA ha558(p1020,p1195,p1200,p1201);
HA ha559(p1197,p1022,p1202,p1203);
HA ha560(p1199,p1201,p1204,p1205);
HA ha561(p1024,p1203,p1206,p1207);
HA ha562(ip_3_15,ip_4_14,p1208,p1209);
HA ha563(ip_5_13,ip_6_12,p1210,p1211);
HA ha564(ip_7_11,ip_8_10,p1212,p1213);
HA ha565(ip_9_9,ip_10_8,p1214,p1215);
HA ha566(ip_11_7,ip_12_6,p1216,p1217);
HA ha567(ip_13_5,ip_14_4,p1218,p1219);
HA ha568(ip_15_3,p1028,p1220,p1221);
HA ha569(p1030,p1032,p1222,p1223);
HA ha570(p1034,p1036,p1224,p1225);
HA ha571(p1209,p1211,p1226,p1227);
HA ha572(p1213,p1215,p1228,p1229);
HA ha573(p1217,p1219,p1230,p1231);
HA ha574(p1038,p1042,p1232,p1233);
HA ha575(p1044,p1046,p1234,p1235);
HA ha576(p1048,p1221,p1236,p1237);
HA ha577(p1223,p1225,p1238,p1239);
HA ha578(p1227,p1229,p1240,p1241);
HA ha579(p1231,p1026,p1242,p1243);
HA ha580(p1050,p1052,p1244,p1245);
HA ha581(p1054,p1056,p1246,p1247);
HA ha582(p1058,p1060,p1248,p1249);
HA ha583(p1233,p1235,p1250,p1251);
HA ha584(p1237,p1239,p1252,p1253);
HA ha585(p1241,p1040,p1254,p1255);
HA ha586(p1062,p1064,p1256,p1257);
HA ha587(p1066,p1068,p1258,p1259);
HA ha588(p1070,p1072,p1260,p1261);
HA ha589(p1243,p1245,p1262,p1263);
HA ha590(p1247,p1249,p1264,p1265);
HA ha591(p1251,p1253,p1266,p1267);
HA ha592(p1074,p1076,p1268,p1269);
HA ha593(p1078,p1080,p1270,p1271);
HA ha594(p1082,p1255,p1272,p1273);
HA ha595(p1257,p1259,p1274,p1275);
HA ha596(p1261,p1263,p1276,p1277);
HA ha597(p1265,p1267,p1278,p1279);
HA ha598(p1084,p1086,p1280,p1281);
HA ha599(p1088,p1090,p1282,p1283);
HA ha600(p1269,p1271,p1284,p1285);
HA ha601(p1273,p1275,p1286,p1287);
HA ha602(p1277,p1279,p1288,p1289);
HA ha603(p1094,p1096,p1290,p1291);
HA ha604(p1098,p1100,p1292,p1293);
HA ha605(p1102,p1281,p1294,p1295);
HA ha606(p1283,p1285,p1296,p1297);
HA ha607(p1287,p1289,p1298,p1299);
HA ha608(p1092,p1104,p1300,p1301);
HA ha609(p1110,p1291,p1302,p1303);
HA ha610(p1293,p1295,p1304,p1305);
HA ha611(p1297,p1299,p1306,p1307);
HA ha612(p1112,p1114,p1308,p1309);
HA ha613(p1116,p1118,p1310,p1311);
HA ha614(p1301,p1303,p1312,p1313);
HA ha615(p1305,p1307,p1314,p1315);
HA ha616(p1106,p1108,p1316,p1317);
HA ha617(p1120,p1122,p1318,p1319);
HA ha618(p1124,p1126,p1320,p1321);
HA ha619(p1128,p1130,p1322,p1323);
HA ha620(p1309,p1311,p1324,p1325);
HA ha621(p1313,p1315,p1326,p1327);
HA ha622(p1132,p1134,p1328,p1329);
HA ha623(p1136,p1138,p1330,p1331);
HA ha624(p1140,p1317,p1332,p1333);
HA ha625(p1319,p1321,p1334,p1335);
HA ha626(p1323,p1325,p1336,p1337);
HA ha627(p1327,p1142,p1338,p1339);
HA ha628(p1144,p1146,p1340,p1341);
HA ha629(p1148,p1150,p1342,p1343);
HA ha630(p1329,p1331,p1344,p1345);
HA ha631(p1333,p1335,p1346,p1347);
HA ha632(p1337,p1152,p1348,p1349);
HA ha633(p1154,p1156,p1350,p1351);
HA ha634(p1158,p1339,p1352,p1353);
FA fa42(p1341,p1343,p1345,p1354,p1355);
HA ha635(p1347,p1160,p1356,p1357);
HA ha636(p1162,p1164,p1358,p1359);
HA ha637(p1166,p1349,p1360,p1361);
HA ha638(p1351,p1353,p1362,p1363);
HA ha639(p1168,p1170,p1364,p1365);
HA ha640(p1172,p1174,p1366,p1367);
HA ha641(p1355,p1357,p1368,p1369);
HA ha642(p1359,p1361,p1370,p1371);
FA fa43(p1363,p1176,p1178,p1372,p1373);
HA ha643(p1180,p1365,p1374,p1375);
HA ha644(p1367,p1369,p1376,p1377);
HA ha645(p1371,p1182,p1378,p1379);
HA ha646(p1184,p1186,p1380,p1381);
HA ha647(p1375,p1377,p1382,p1383);
HA ha648(p1190,p1373,p1384,p1385);
HA ha649(p1379,p1381,p1386,p1387);
HA ha650(p1383,p1192,p1388,p1389);
HA ha651(p1385,p1387,p1390,p1391);
HA ha652(p1188,p1194,p1392,p1393);
HA ha653(p1196,p1389,p1394,p1395);
HA ha654(p1391,p1198,p1396,p1397);
FA fa44(p1200,p1393,p1395,p1398,p1399);
HA ha655(p1202,p1204,p1400,p1401);
HA ha656(p1397,p1206,p1402,p1403);
HA ha657(p1399,p1401,p1404,p1405);
HA ha658(ip_4_15,ip_5_14,p1406,p1407);
HA ha659(ip_6_13,ip_7_12,p1408,p1409);
HA ha660(ip_8_11,ip_9_10,p1410,p1411);
HA ha661(ip_10_9,ip_11_8,p1412,p1413);
HA ha662(ip_12_7,ip_13_6,p1414,p1415);
HA ha663(ip_14_5,ip_15_4,p1416,p1417);
HA ha664(p1208,p1210,p1418,p1419);
HA ha665(p1212,p1214,p1420,p1421);
HA ha666(p1216,p1218,p1422,p1423);
HA ha667(p1407,p1409,p1424,p1425);
HA ha668(p1411,p1413,p1426,p1427);
HA ha669(p1415,p1417,p1428,p1429);
HA ha670(p1220,p1222,p1430,p1431);
HA ha671(p1224,p1226,p1432,p1433);
HA ha672(p1228,p1230,p1434,p1435);
HA ha673(p1419,p1421,p1436,p1437);
HA ha674(p1423,p1425,p1438,p1439);
HA ha675(p1427,p1429,p1440,p1441);
HA ha676(p1232,p1234,p1442,p1443);
HA ha677(p1236,p1238,p1444,p1445);
HA ha678(p1240,p1431,p1446,p1447);
HA ha679(p1433,p1435,p1448,p1449);
HA ha680(p1437,p1439,p1450,p1451);
FA fa45(p1441,p1242,p1244,p1452,p1453);
HA ha681(p1246,p1248,p1454,p1455);
HA ha682(p1250,p1252,p1456,p1457);
HA ha683(p1443,p1445,p1458,p1459);
FA fa46(p1447,p1449,p1451,p1460,p1461);
HA ha684(p1254,p1256,p1462,p1463);
HA ha685(p1258,p1260,p1464,p1465);
HA ha686(p1262,p1264,p1466,p1467);
HA ha687(p1266,p1455,p1468,p1469);
HA ha688(p1457,p1459,p1470,p1471);
HA ha689(p1268,p1270,p1472,p1473);
HA ha690(p1272,p1274,p1474,p1475);
HA ha691(p1276,p1278,p1476,p1477);
HA ha692(p1453,p1461,p1478,p1479);
HA ha693(p1463,p1465,p1480,p1481);
HA ha694(p1467,p1469,p1482,p1483);
HA ha695(p1471,p1280,p1484,p1485);
HA ha696(p1282,p1284,p1486,p1487);
HA ha697(p1286,p1288,p1488,p1489);
HA ha698(p1473,p1475,p1490,p1491);
HA ha699(p1477,p1479,p1492,p1493);
HA ha700(p1481,p1483,p1494,p1495);
HA ha701(p1290,p1292,p1496,p1497);
FA fa47(p1294,p1296,p1298,p1498,p1499);
HA ha702(p1485,p1487,p1500,p1501);
HA ha703(p1489,p1491,p1502,p1503);
HA ha704(p1493,p1495,p1504,p1505);
HA ha705(p1300,p1302,p1506,p1507);
HA ha706(p1304,p1306,p1508,p1509);
HA ha707(p1497,p1501,p1510,p1511);
FA fa48(p1503,p1505,p1308,p1512,p1513);
HA ha708(p1310,p1312,p1514,p1515);
HA ha709(p1314,p1499,p1516,p1517);
HA ha710(p1507,p1509,p1518,p1519);
HA ha711(p1511,p1316,p1520,p1521);
HA ha712(p1318,p1320,p1522,p1523);
HA ha713(p1322,p1324,p1524,p1525);
HA ha714(p1326,p1513,p1526,p1527);
HA ha715(p1515,p1517,p1528,p1529);
HA ha716(p1519,p1328,p1530,p1531);
HA ha717(p1330,p1332,p1532,p1533);
FA fa49(p1334,p1336,p1521,p1534,p1535);
HA ha718(p1523,p1525,p1536,p1537);
HA ha719(p1527,p1529,p1538,p1539);
HA ha720(p1338,p1340,p1540,p1541);
HA ha721(p1342,p1344,p1542,p1543);
HA ha722(p1346,p1531,p1544,p1545);
HA ha723(p1533,p1537,p1546,p1547);
HA ha724(p1539,p1348,p1548,p1549);
HA ha725(p1350,p1352,p1550,p1551);
HA ha726(p1535,p1541,p1552,p1553);
HA ha727(p1543,p1545,p1554,p1555);
HA ha728(p1547,p1356,p1556,p1557);
FA fa50(p1358,p1360,p1362,p1558,p1559);
HA ha729(p1549,p1551,p1560,p1561);
HA ha730(p1553,p1555,p1562,p1563);
HA ha731(p1354,p1364,p1564,p1565);
HA ha732(p1366,p1368,p1566,p1567);
HA ha733(p1370,p1557,p1568,p1569);
HA ha734(p1561,p1563,p1570,p1571);
HA ha735(p1374,p1376,p1572,p1573);
HA ha736(p1559,p1565,p1574,p1575);
HA ha737(p1567,p1569,p1576,p1577);
HA ha738(p1571,p1378,p1578,p1579);
HA ha739(p1380,p1382,p1580,p1581);
HA ha740(p1573,p1575,p1582,p1583);
HA ha741(p1577,p1372,p1584,p1585);
HA ha742(p1384,p1386,p1586,p1587);
HA ha743(p1579,p1581,p1588,p1589);
HA ha744(p1583,p1388,p1590,p1591);
HA ha745(p1390,p1585,p1592,p1593);
HA ha746(p1587,p1589,p1594,p1595);
HA ha747(p1392,p1394,p1596,p1597);
HA ha748(p1591,p1593,p1598,p1599);
HA ha749(p1595,p1396,p1600,p1601);
HA ha750(p1597,p1599,p1602,p1603);
HA ha751(p1400,p1601,p1604,p1605);
HA ha752(p1603,p1398,p1606,p1607);
HA ha753(p1402,p1404,p1608,p1609);
HA ha754(p1605,p1607,p1610,p1611);
HA ha755(ip_5_15,ip_6_14,p1612,p1613);
FA fa51(ip_7_13,ip_8_12,ip_9_11,p1614,p1615);
FA fa52(ip_10_10,ip_11_9,ip_12_8,p1616,p1617);
HA ha756(ip_13_7,ip_14_6,p1618,p1619);
FA fa53(ip_15_5,p1406,p1408,p1620,p1621);
HA ha757(p1410,p1412,p1622,p1623);
HA ha758(p1414,p1416,p1624,p1625);
HA ha759(p1613,p1619,p1626,p1627);
HA ha760(p1418,p1420,p1628,p1629);
HA ha761(p1422,p1424,p1630,p1631);
HA ha762(p1426,p1428,p1632,p1633);
HA ha763(p1615,p1617,p1634,p1635);
HA ha764(p1623,p1625,p1636,p1637);
HA ha765(p1627,p1430,p1638,p1639);
HA ha766(p1432,p1434,p1640,p1641);
HA ha767(p1436,p1438,p1642,p1643);
HA ha768(p1440,p1621,p1644,p1645);
HA ha769(p1629,p1631,p1646,p1647);
FA fa54(p1633,p1635,p1637,p1648,p1649);
HA ha770(p1442,p1444,p1650,p1651);
HA ha771(p1446,p1448,p1652,p1653);
HA ha772(p1450,p1639,p1654,p1655);
HA ha773(p1641,p1643,p1656,p1657);
HA ha774(p1645,p1647,p1658,p1659);
HA ha775(p1454,p1456,p1660,p1661);
HA ha776(p1458,p1649,p1662,p1663);
HA ha777(p1651,p1653,p1664,p1665);
HA ha778(p1655,p1657,p1666,p1667);
HA ha779(p1659,p1462,p1668,p1669);
HA ha780(p1464,p1466,p1670,p1671);
HA ha781(p1468,p1470,p1672,p1673);
HA ha782(p1661,p1663,p1674,p1675);
HA ha783(p1665,p1667,p1676,p1677);
HA ha784(p1452,p1460,p1678,p1679);
HA ha785(p1472,p1474,p1680,p1681);
HA ha786(p1476,p1478,p1682,p1683);
HA ha787(p1480,p1482,p1684,p1685);
HA ha788(p1669,p1671,p1686,p1687);
HA ha789(p1673,p1675,p1688,p1689);
HA ha790(p1677,p1484,p1690,p1691);
HA ha791(p1486,p1488,p1692,p1693);
HA ha792(p1490,p1492,p1694,p1695);
HA ha793(p1494,p1679,p1696,p1697);
HA ha794(p1681,p1683,p1698,p1699);
HA ha795(p1685,p1687,p1700,p1701);
HA ha796(p1689,p1496,p1702,p1703);
HA ha797(p1500,p1502,p1704,p1705);
HA ha798(p1504,p1691,p1706,p1707);
HA ha799(p1693,p1695,p1708,p1709);
HA ha800(p1697,p1699,p1710,p1711);
HA ha801(p1701,p1506,p1712,p1713);
HA ha802(p1508,p1510,p1714,p1715);
HA ha803(p1703,p1705,p1716,p1717);
HA ha804(p1707,p1709,p1718,p1719);
HA ha805(p1711,p1498,p1720,p1721);
HA ha806(p1514,p1516,p1722,p1723);
HA ha807(p1518,p1713,p1724,p1725);
HA ha808(p1715,p1717,p1726,p1727);
HA ha809(p1719,p1512,p1728,p1729);
HA ha810(p1520,p1522,p1730,p1731);
HA ha811(p1524,p1526,p1732,p1733);
HA ha812(p1528,p1721,p1734,p1735);
HA ha813(p1723,p1725,p1736,p1737);
HA ha814(p1727,p1530,p1738,p1739);
FA fa55(p1532,p1536,p1538,p1740,p1741);
HA ha815(p1729,p1731,p1742,p1743);
HA ha816(p1733,p1735,p1744,p1745);
HA ha817(p1737,p1540,p1746,p1747);
HA ha818(p1542,p1544,p1748,p1749);
HA ha819(p1546,p1739,p1750,p1751);
HA ha820(p1743,p1745,p1752,p1753);
HA ha821(p1534,p1548,p1754,p1755);
HA ha822(p1550,p1552,p1756,p1757);
HA ha823(p1554,p1741,p1758,p1759);
HA ha824(p1747,p1749,p1760,p1761);
HA ha825(p1751,p1753,p1762,p1763);
HA ha826(p1556,p1560,p1764,p1765);
HA ha827(p1562,p1755,p1766,p1767);
HA ha828(p1757,p1759,p1768,p1769);
HA ha829(p1761,p1763,p1770,p1771);
HA ha830(p1564,p1566,p1772,p1773);
HA ha831(p1568,p1570,p1774,p1775);
HA ha832(p1765,p1767,p1776,p1777);
HA ha833(p1769,p1771,p1778,p1779);
HA ha834(p1558,p1572,p1780,p1781);
HA ha835(p1574,p1576,p1782,p1783);
HA ha836(p1773,p1775,p1784,p1785);
HA ha837(p1777,p1779,p1786,p1787);
HA ha838(p1578,p1580,p1788,p1789);
HA ha839(p1582,p1781,p1790,p1791);
HA ha840(p1783,p1785,p1792,p1793);
HA ha841(p1787,p1584,p1794,p1795);
HA ha842(p1586,p1588,p1796,p1797);
HA ha843(p1789,p1791,p1798,p1799);
HA ha844(p1793,p1590,p1800,p1801);
HA ha845(p1592,p1594,p1802,p1803);
HA ha846(p1795,p1797,p1804,p1805);
HA ha847(p1799,p1596,p1806,p1807);
HA ha848(p1598,p1801,p1808,p1809);
HA ha849(p1803,p1805,p1810,p1811);
HA ha850(p1600,p1602,p1812,p1813);
HA ha851(p1807,p1809,p1814,p1815);
HA ha852(p1811,p1604,p1816,p1817);
HA ha853(p1813,p1815,p1818,p1819);
HA ha854(p1606,p1608,p1820,p1821);
HA ha855(p1817,p1819,p1822,p1823);
HA ha856(p1610,p1821,p1824,p1825);
HA ha857(ip_6_15,ip_7_14,p1826,p1827);
HA ha858(ip_8_13,ip_9_12,p1828,p1829);
HA ha859(ip_10_11,ip_11_10,p1830,p1831);
HA ha860(ip_12_9,ip_13_8,p1832,p1833);
HA ha861(ip_14_7,ip_15_6,p1834,p1835);
HA ha862(p1612,p1618,p1836,p1837);
HA ha863(p1827,p1829,p1838,p1839);
HA ha864(p1831,p1833,p1840,p1841);
HA ha865(p1835,p1622,p1842,p1843);
HA ha866(p1624,p1626,p1844,p1845);
HA ha867(p1837,p1839,p1846,p1847);
HA ha868(p1841,p1614,p1848,p1849);
HA ha869(p1616,p1628,p1850,p1851);
HA ha870(p1630,p1632,p1852,p1853);
HA ha871(p1634,p1636,p1854,p1855);
HA ha872(p1843,p1845,p1856,p1857);
HA ha873(p1847,p1620,p1858,p1859);
HA ha874(p1638,p1640,p1860,p1861);
HA ha875(p1642,p1644,p1862,p1863);
HA ha876(p1646,p1849,p1864,p1865);
HA ha877(p1851,p1853,p1866,p1867);
HA ha878(p1855,p1857,p1868,p1869);
HA ha879(p1650,p1652,p1870,p1871);
HA ha880(p1654,p1656,p1872,p1873);
HA ha881(p1658,p1859,p1874,p1875);
HA ha882(p1861,p1863,p1876,p1877);
HA ha883(p1865,p1867,p1878,p1879);
FA fa56(p1869,p1648,p1660,p1880,p1881);
HA ha884(p1662,p1664,p1882,p1883);
HA ha885(p1666,p1871,p1884,p1885);
HA ha886(p1873,p1875,p1886,p1887);
HA ha887(p1877,p1879,p1888,p1889);
HA ha888(p1668,p1670,p1890,p1891);
HA ha889(p1672,p1674,p1892,p1893);
HA ha890(p1676,p1883,p1894,p1895);
HA ha891(p1885,p1887,p1896,p1897);
HA ha892(p1889,p1678,p1898,p1899);
HA ha893(p1680,p1682,p1900,p1901);
HA ha894(p1684,p1686,p1902,p1903);
HA ha895(p1688,p1881,p1904,p1905);
HA ha896(p1891,p1893,p1906,p1907);
HA ha897(p1895,p1897,p1908,p1909);
HA ha898(p1690,p1692,p1910,p1911);
HA ha899(p1694,p1696,p1912,p1913);
HA ha900(p1698,p1700,p1914,p1915);
HA ha901(p1899,p1901,p1916,p1917);
HA ha902(p1903,p1905,p1918,p1919);
HA ha903(p1907,p1909,p1920,p1921);
HA ha904(p1702,p1704,p1922,p1923);
HA ha905(p1706,p1708,p1924,p1925);
FA fa57(p1710,p1911,p1913,p1926,p1927);
HA ha906(p1915,p1917,p1928,p1929);
HA ha907(p1919,p1921,p1930,p1931);
HA ha908(p1712,p1714,p1932,p1933);
HA ha909(p1716,p1718,p1934,p1935);
HA ha910(p1923,p1925,p1936,p1937);
HA ha911(p1929,p1931,p1938,p1939);
HA ha912(p1720,p1722,p1940,p1941);
HA ha913(p1724,p1726,p1942,p1943);
HA ha914(p1927,p1933,p1944,p1945);
HA ha915(p1935,p1937,p1946,p1947);
HA ha916(p1939,p1728,p1948,p1949);
FA fa58(p1730,p1732,p1734,p1950,p1951);
HA ha917(p1736,p1941,p1952,p1953);
FA fa59(p1943,p1945,p1947,p1954,p1955);
HA ha918(p1738,p1742,p1956,p1957);
HA ha919(p1744,p1949,p1958,p1959);
HA ha920(p1953,p1746,p1960,p1961);
HA ha921(p1748,p1750,p1962,p1963);
HA ha922(p1752,p1951,p1964,p1965);
HA ha923(p1955,p1957,p1966,p1967);
HA ha924(p1959,p1740,p1968,p1969);
HA ha925(p1754,p1756,p1970,p1971);
HA ha926(p1758,p1760,p1972,p1973);
HA ha927(p1762,p1961,p1974,p1975);
HA ha928(p1963,p1965,p1976,p1977);
HA ha929(p1967,p1764,p1978,p1979);
HA ha930(p1766,p1768,p1980,p1981);
HA ha931(p1770,p1969,p1982,p1983);
HA ha932(p1971,p1973,p1984,p1985);
HA ha933(p1975,p1977,p1986,p1987);
HA ha934(p1772,p1774,p1988,p1989);
HA ha935(p1776,p1778,p1990,p1991);
HA ha936(p1979,p1981,p1992,p1993);
HA ha937(p1983,p1985,p1994,p1995);
HA ha938(p1987,p1780,p1996,p1997);
HA ha939(p1782,p1784,p1998,p1999);
HA ha940(p1786,p1989,p2000,p2001);
HA ha941(p1991,p1993,p2002,p2003);
HA ha942(p1995,p1788,p2004,p2005);
HA ha943(p1790,p1792,p2006,p2007);
HA ha944(p1997,p1999,p2008,p2009);
HA ha945(p2001,p2003,p2010,p2011);
HA ha946(p1794,p1796,p2012,p2013);
HA ha947(p1798,p2005,p2014,p2015);
HA ha948(p2007,p2009,p2016,p2017);
HA ha949(p2011,p1800,p2018,p2019);
HA ha950(p1802,p1804,p2020,p2021);
HA ha951(p2013,p2015,p2022,p2023);
FA fa60(p2017,p1806,p1808,p2024,p2025);
HA ha952(p1810,p2019,p2026,p2027);
HA ha953(p2021,p2023,p2028,p2029);
HA ha954(p1812,p1814,p2030,p2031);
HA ha955(p2027,p2029,p2032,p2033);
HA ha956(p1816,p1818,p2034,p2035);
HA ha957(p2025,p2031,p2036,p2037);
HA ha958(p2033,p1820,p2038,p2039);
HA ha959(p1822,p2035,p2040,p2041);
HA ha960(p2037,p1824,p2042,p2043);
HA ha961(p2039,p2041,p2044,p2045);
HA ha962(ip_7_15,ip_8_14,p2046,p2047);
HA ha963(ip_9_13,ip_10_12,p2048,p2049);
HA ha964(ip_11_11,ip_12_10,p2050,p2051);
HA ha965(ip_13_9,ip_14_8,p2052,p2053);
HA ha966(ip_15_7,p1826,p2054,p2055);
HA ha967(p1828,p1830,p2056,p2057);
HA ha968(p1832,p1834,p2058,p2059);
HA ha969(p2047,p2049,p2060,p2061);
HA ha970(p2051,p2053,p2062,p2063);
HA ha971(p1836,p1838,p2064,p2065);
HA ha972(p1840,p2055,p2066,p2067);
HA ha973(p2057,p2059,p2068,p2069);
HA ha974(p2061,p2063,p2070,p2071);
HA ha975(p1842,p1844,p2072,p2073);
HA ha976(p1846,p2065,p2074,p2075);
HA ha977(p2067,p2069,p2076,p2077);
HA ha978(p2071,p1848,p2078,p2079);
HA ha979(p1850,p1852,p2080,p2081);
HA ha980(p1854,p1856,p2082,p2083);
HA ha981(p2073,p2075,p2084,p2085);
HA ha982(p2077,p1858,p2086,p2087);
HA ha983(p1860,p1862,p2088,p2089);
HA ha984(p1864,p1866,p2090,p2091);
FA fa61(p1868,p2079,p2081,p2092,p2093);
HA ha985(p2083,p2085,p2094,p2095);
HA ha986(p1870,p1872,p2096,p2097);
HA ha987(p1874,p1876,p2098,p2099);
HA ha988(p1878,p2087,p2100,p2101);
HA ha989(p2089,p2091,p2102,p2103);
HA ha990(p2095,p1882,p2104,p2105);
HA ha991(p1884,p1886,p2106,p2107);
FA fa62(p1888,p2093,p2097,p2108,p2109);
HA ha992(p2099,p2101,p2110,p2111);
HA ha993(p2103,p1890,p2112,p2113);
HA ha994(p1892,p1894,p2114,p2115);
HA ha995(p1896,p2105,p2116,p2117);
HA ha996(p2107,p2111,p2118,p2119);
HA ha997(p1880,p1898,p2120,p2121);
HA ha998(p1900,p1902,p2122,p2123);
HA ha999(p1904,p1906,p2124,p2125);
HA ha1000(p1908,p2109,p2126,p2127);
HA ha1001(p2113,p2115,p2128,p2129);
HA ha1002(p2117,p2119,p2130,p2131);
HA ha1003(p1910,p1912,p2132,p2133);
HA ha1004(p1914,p1916,p2134,p2135);
HA ha1005(p1918,p1920,p2136,p2137);
HA ha1006(p2121,p2123,p2138,p2139);
HA ha1007(p2125,p2127,p2140,p2141);
HA ha1008(p2129,p2131,p2142,p2143);
HA ha1009(p1922,p1924,p2144,p2145);
HA ha1010(p1928,p1930,p2146,p2147);
HA ha1011(p2133,p2135,p2148,p2149);
HA ha1012(p2137,p2139,p2150,p2151);
HA ha1013(p2141,p2143,p2152,p2153);
HA ha1014(p1932,p1934,p2154,p2155);
HA ha1015(p1936,p1938,p2156,p2157);
HA ha1016(p2145,p2147,p2158,p2159);
HA ha1017(p2149,p2151,p2160,p2161);
HA ha1018(p2153,p1926,p2162,p2163);
HA ha1019(p1940,p1942,p2164,p2165);
HA ha1020(p1944,p1946,p2166,p2167);
HA ha1021(p2155,p2157,p2168,p2169);
HA ha1022(p2159,p2161,p2170,p2171);
HA ha1023(p1948,p1952,p2172,p2173);
HA ha1024(p2163,p2165,p2174,p2175);
HA ha1025(p2167,p2169,p2176,p2177);
HA ha1026(p2171,p1956,p2178,p2179);
HA ha1027(p1958,p2173,p2180,p2181);
HA ha1028(p2175,p2177,p2182,p2183);
HA ha1029(p1950,p1954,p2184,p2185);
HA ha1030(p1960,p1962,p2186,p2187);
FA fa63(p1964,p1966,p2179,p2188,p2189);
HA ha1031(p2181,p2183,p2190,p2191);
HA ha1032(p1968,p1970,p2192,p2193);
HA ha1033(p1972,p1974,p2194,p2195);
HA ha1034(p1976,p2185,p2196,p2197);
HA ha1035(p2187,p2191,p2198,p2199);
HA ha1036(p1978,p1980,p2200,p2201);
HA ha1037(p1982,p1984,p2202,p2203);
HA ha1038(p1986,p2189,p2204,p2205);
HA ha1039(p2193,p2195,p2206,p2207);
HA ha1040(p2197,p2199,p2208,p2209);
HA ha1041(p1988,p1990,p2210,p2211);
HA ha1042(p1992,p1994,p2212,p2213);
HA ha1043(p2201,p2203,p2214,p2215);
HA ha1044(p2205,p2207,p2216,p2217);
HA ha1045(p2209,p1996,p2218,p2219);
HA ha1046(p1998,p2000,p2220,p2221);
HA ha1047(p2002,p2211,p2222,p2223);
HA ha1048(p2213,p2215,p2224,p2225);
HA ha1049(p2217,p2004,p2226,p2227);
HA ha1050(p2006,p2008,p2228,p2229);
HA ha1051(p2010,p2219,p2230,p2231);
HA ha1052(p2221,p2223,p2232,p2233);
HA ha1053(p2225,p2012,p2234,p2235);
FA fa64(p2014,p2016,p2227,p2236,p2237);
HA ha1054(p2229,p2231,p2238,p2239);
HA ha1055(p2233,p2018,p2240,p2241);
HA ha1056(p2020,p2022,p2242,p2243);
HA ha1057(p2235,p2239,p2244,p2245);
HA ha1058(p2026,p2028,p2246,p2247);
HA ha1059(p2237,p2241,p2248,p2249);
HA ha1060(p2243,p2245,p2250,p2251);
HA ha1061(p2030,p2032,p2252,p2253);
HA ha1062(p2247,p2249,p2254,p2255);
HA ha1063(p2251,p2024,p2256,p2257);
HA ha1064(p2034,p2036,p2258,p2259);
HA ha1065(p2253,p2255,p2260,p2261);
HA ha1066(p2038,p2040,p2262,p2263);
HA ha1067(p2257,p2259,p2264,p2265);
HA ha1068(p2261,p2042,p2266,p2267);
HA ha1069(p2044,p2263,p2268,p2269);
HA ha1070(p2265,p2267,p2270,p2271);
HA ha1071(ip_8_15,ip_9_14,p2272,p2273);
HA ha1072(ip_10_13,ip_11_12,p2274,p2275);
HA ha1073(ip_12_11,ip_13_10,p2276,p2277);
HA ha1074(ip_14_9,ip_15_8,p2278,p2279);
FA fa65(p2046,p2048,p2050,p2280,p2281);
HA ha1075(p2052,p2273,p2282,p2283);
HA ha1076(p2275,p2277,p2284,p2285);
HA ha1077(p2279,p2054,p2286,p2287);
HA ha1078(p2056,p2058,p2288,p2289);
HA ha1079(p2060,p2062,p2290,p2291);
HA ha1080(p2283,p2285,p2292,p2293);
FA fa66(p2064,p2066,p2068,p2294,p2295);
HA ha1081(p2070,p2281,p2296,p2297);
HA ha1082(p2287,p2289,p2298,p2299);
HA ha1083(p2291,p2293,p2300,p2301);
HA ha1084(p2072,p2074,p2302,p2303);
HA ha1085(p2076,p2297,p2304,p2305);
HA ha1086(p2299,p2301,p2306,p2307);
HA ha1087(p2078,p2080,p2308,p2309);
HA ha1088(p2082,p2084,p2310,p2311);
HA ha1089(p2295,p2303,p2312,p2313);
HA ha1090(p2305,p2307,p2314,p2315);
HA ha1091(p2086,p2088,p2316,p2317);
HA ha1092(p2090,p2094,p2318,p2319);
HA ha1093(p2309,p2311,p2320,p2321);
HA ha1094(p2313,p2315,p2322,p2323);
HA ha1095(p2096,p2098,p2324,p2325);
HA ha1096(p2100,p2102,p2326,p2327);
HA ha1097(p2317,p2319,p2328,p2329);
HA ha1098(p2321,p2323,p2330,p2331);
HA ha1099(p2092,p2104,p2332,p2333);
HA ha1100(p2106,p2110,p2334,p2335);
HA ha1101(p2325,p2327,p2336,p2337);
HA ha1102(p2329,p2331,p2338,p2339);
FA fa67(p2112,p2114,p2116,p2340,p2341);
HA ha1103(p2118,p2333,p2342,p2343);
HA ha1104(p2335,p2337,p2344,p2345);
HA ha1105(p2339,p2108,p2346,p2347);
HA ha1106(p2120,p2122,p2348,p2349);
HA ha1107(p2124,p2126,p2350,p2351);
HA ha1108(p2128,p2130,p2352,p2353);
HA ha1109(p2343,p2345,p2354,p2355);
HA ha1110(p2132,p2134,p2356,p2357);
HA ha1111(p2136,p2138,p2358,p2359);
HA ha1112(p2140,p2142,p2360,p2361);
HA ha1113(p2341,p2347,p2362,p2363);
HA ha1114(p2349,p2351,p2364,p2365);
HA ha1115(p2353,p2355,p2366,p2367);
HA ha1116(p2144,p2146,p2368,p2369);
HA ha1117(p2148,p2150,p2370,p2371);
HA ha1118(p2152,p2357,p2372,p2373);
HA ha1119(p2359,p2361,p2374,p2375);
HA ha1120(p2363,p2365,p2376,p2377);
HA ha1121(p2367,p2154,p2378,p2379);
HA ha1122(p2156,p2158,p2380,p2381);
HA ha1123(p2160,p2369,p2382,p2383);
HA ha1124(p2371,p2373,p2384,p2385);
FA fa68(p2375,p2377,p2162,p2386,p2387);
HA ha1125(p2164,p2166,p2388,p2389);
FA fa69(p2168,p2170,p2379,p2390,p2391);
HA ha1126(p2381,p2383,p2392,p2393);
HA ha1127(p2385,p2172,p2394,p2395);
HA ha1128(p2174,p2176,p2396,p2397);
HA ha1129(p2387,p2389,p2398,p2399);
HA ha1130(p2393,p2178,p2400,p2401);
HA ha1131(p2180,p2182,p2402,p2403);
HA ha1132(p2391,p2395,p2404,p2405);
HA ha1133(p2397,p2399,p2406,p2407);
HA ha1134(p2184,p2186,p2408,p2409);
HA ha1135(p2190,p2401,p2410,p2411);
HA ha1136(p2403,p2405,p2412,p2413);
HA ha1137(p2407,p2192,p2414,p2415);
HA ha1138(p2194,p2196,p2416,p2417);
HA ha1139(p2198,p2409,p2418,p2419);
FA fa70(p2411,p2413,p2188,p2420,p2421);
HA ha1140(p2200,p2202,p2422,p2423);
HA ha1141(p2204,p2206,p2424,p2425);
FA fa71(p2208,p2415,p2417,p2426,p2427);
HA ha1142(p2419,p2210,p2428,p2429);
FA fa72(p2212,p2214,p2216,p2430,p2431);
HA ha1143(p2421,p2423,p2432,p2433);
HA ha1144(p2425,p2218,p2434,p2435);
FA fa73(p2220,p2222,p2224,p2436,p2437);
HA ha1145(p2427,p2429,p2438,p2439);
HA ha1146(p2433,p2226,p2440,p2441);
HA ha1147(p2228,p2230,p2442,p2443);
HA ha1148(p2232,p2431,p2444,p2445);
HA ha1149(p2435,p2439,p2446,p2447);
HA ha1150(p2234,p2238,p2448,p2449);
HA ha1151(p2437,p2441,p2450,p2451);
HA ha1152(p2443,p2445,p2452,p2453);
HA ha1153(p2447,p2240,p2454,p2455);
HA ha1154(p2242,p2244,p2456,p2457);
HA ha1155(p2449,p2451,p2458,p2459);
HA ha1156(p2453,p2236,p2460,p2461);
HA ha1157(p2246,p2248,p2462,p2463);
HA ha1158(p2250,p2455,p2464,p2465);
HA ha1159(p2457,p2459,p2466,p2467);
HA ha1160(p2252,p2254,p2468,p2469);
HA ha1161(p2461,p2463,p2470,p2471);
HA ha1162(p2465,p2467,p2472,p2473);
HA ha1163(p2256,p2258,p2474,p2475);
HA ha1164(p2260,p2469,p2476,p2477);
HA ha1165(p2471,p2473,p2478,p2479);
HA ha1166(p2262,p2264,p2480,p2481);
HA ha1167(p2475,p2477,p2482,p2483);
HA ha1168(p2479,p2266,p2484,p2485);
HA ha1169(p2268,p2481,p2486,p2487);
HA ha1170(p2483,p2270,p2488,p2489);
HA ha1171(p2485,p2487,p2490,p2491);
HA ha1172(ip_9_15,ip_10_14,p2492,p2493);
FA fa74(ip_11_13,ip_12_12,ip_13_11,p2494,p2495);
HA ha1173(ip_14_10,ip_15_9,p2496,p2497);
HA ha1174(p2272,p2274,p2498,p2499);
HA ha1175(p2276,p2278,p2500,p2501);
HA ha1176(p2493,p2497,p2502,p2503);
HA ha1177(p2282,p2284,p2504,p2505);
HA ha1178(p2495,p2499,p2506,p2507);
HA ha1179(p2501,p2503,p2508,p2509);
HA ha1180(p2286,p2288,p2510,p2511);
FA fa75(p2290,p2292,p2505,p2512,p2513);
HA ha1181(p2507,p2509,p2514,p2515);
HA ha1182(p2280,p2296,p2516,p2517);
HA ha1183(p2298,p2300,p2518,p2519);
HA ha1184(p2511,p2515,p2520,p2521);
HA ha1185(p2302,p2304,p2522,p2523);
HA ha1186(p2306,p2513,p2524,p2525);
HA ha1187(p2517,p2519,p2526,p2527);
HA ha1188(p2521,p2294,p2528,p2529);
HA ha1189(p2308,p2310,p2530,p2531);
HA ha1190(p2312,p2314,p2532,p2533);
HA ha1191(p2523,p2525,p2534,p2535);
HA ha1192(p2527,p2316,p2536,p2537);
HA ha1193(p2318,p2320,p2538,p2539);
HA ha1194(p2322,p2529,p2540,p2541);
HA ha1195(p2531,p2533,p2542,p2543);
HA ha1196(p2535,p2324,p2544,p2545);
HA ha1197(p2326,p2328,p2546,p2547);
HA ha1198(p2330,p2537,p2548,p2549);
FA fa76(p2539,p2541,p2543,p2550,p2551);
HA ha1199(p2332,p2334,p2552,p2553);
HA ha1200(p2336,p2338,p2554,p2555);
HA ha1201(p2545,p2547,p2556,p2557);
HA ha1202(p2549,p2342,p2558,p2559);
HA ha1203(p2344,p2551,p2560,p2561);
HA ha1204(p2553,p2555,p2562,p2563);
HA ha1205(p2557,p2346,p2564,p2565);
HA ha1206(p2348,p2350,p2566,p2567);
HA ha1207(p2352,p2354,p2568,p2569);
HA ha1208(p2559,p2561,p2570,p2571);
FA fa77(p2563,p2340,p2356,p2572,p2573);
HA ha1209(p2358,p2360,p2574,p2575);
HA ha1210(p2362,p2364,p2576,p2577);
HA ha1211(p2366,p2565,p2578,p2579);
HA ha1212(p2567,p2569,p2580,p2581);
HA ha1213(p2571,p2368,p2582,p2583);
HA ha1214(p2370,p2372,p2584,p2585);
HA ha1215(p2374,p2376,p2586,p2587);
HA ha1216(p2575,p2577,p2588,p2589);
HA ha1217(p2579,p2581,p2590,p2591);
HA ha1218(p2378,p2380,p2592,p2593);
HA ha1219(p2382,p2384,p2594,p2595);
HA ha1220(p2573,p2583,p2596,p2597);
HA ha1221(p2585,p2587,p2598,p2599);
FA fa78(p2589,p2591,p2388,p2600,p2601);
HA ha1222(p2392,p2593,p2602,p2603);
HA ha1223(p2595,p2597,p2604,p2605);
HA ha1224(p2599,p2386,p2606,p2607);
HA ha1225(p2394,p2396,p2608,p2609);
HA ha1226(p2398,p2601,p2610,p2611);
HA ha1227(p2603,p2605,p2612,p2613);
HA ha1228(p2390,p2400,p2614,p2615);
HA ha1229(p2402,p2404,p2616,p2617);
HA ha1230(p2406,p2607,p2618,p2619);
FA fa79(p2609,p2611,p2613,p2620,p2621);
FA fa80(p2408,p2410,p2412,p2622,p2623);
HA ha1231(p2615,p2617,p2624,p2625);
HA ha1232(p2619,p2414,p2626,p2627);
HA ha1233(p2416,p2418,p2628,p2629);
HA ha1234(p2621,p2625,p2630,p2631);
HA ha1235(p2422,p2424,p2632,p2633);
HA ha1236(p2623,p2627,p2634,p2635);
HA ha1237(p2629,p2631,p2636,p2637);
HA ha1238(p2420,p2428,p2638,p2639);
HA ha1239(p2432,p2633,p2640,p2641);
HA ha1240(p2635,p2637,p2642,p2643);
HA ha1241(p2426,p2434,p2644,p2645);
HA ha1242(p2438,p2639,p2646,p2647);
HA ha1243(p2641,p2643,p2648,p2649);
HA ha1244(p2430,p2440,p2650,p2651);
HA ha1245(p2442,p2444,p2652,p2653);
HA ha1246(p2446,p2645,p2654,p2655);
HA ha1247(p2647,p2649,p2656,p2657);
HA ha1248(p2436,p2448,p2658,p2659);
HA ha1249(p2450,p2452,p2660,p2661);
HA ha1250(p2651,p2653,p2662,p2663);
HA ha1251(p2655,p2657,p2664,p2665);
HA ha1252(p2454,p2456,p2666,p2667);
FA fa81(p2458,p2659,p2661,p2668,p2669);
HA ha1253(p2663,p2665,p2670,p2671);
HA ha1254(p2460,p2462,p2672,p2673);
HA ha1255(p2464,p2466,p2674,p2675);
HA ha1256(p2667,p2671,p2676,p2677);
HA ha1257(p2468,p2470,p2678,p2679);
HA ha1258(p2472,p2669,p2680,p2681);
HA ha1259(p2673,p2675,p2682,p2683);
HA ha1260(p2677,p2474,p2684,p2685);
HA ha1261(p2476,p2478,p2686,p2687);
HA ha1262(p2679,p2681,p2688,p2689);
HA ha1263(p2683,p2480,p2690,p2691);
HA ha1264(p2482,p2685,p2692,p2693);
HA ha1265(p2687,p2689,p2694,p2695);
HA ha1266(p2484,p2486,p2696,p2697);
HA ha1267(p2691,p2693,p2698,p2699);
HA ha1268(p2695,p2488,p2700,p2701);
HA ha1269(p2490,p2697,p2702,p2703);
HA ha1270(p2699,p2701,p2704,p2705);
HA ha1271(ip_10_15,ip_11_14,p2706,p2707);
HA ha1272(ip_12_13,ip_13_12,p2708,p2709);
HA ha1273(ip_14_11,ip_15_10,p2710,p2711);
HA ha1274(p2492,p2496,p2712,p2713);
HA ha1275(p2707,p2709,p2714,p2715);
HA ha1276(p2711,p2498,p2716,p2717);
FA fa82(p2500,p2502,p2713,p2718,p2719);
HA ha1277(p2715,p2494,p2720,p2721);
FA fa83(p2504,p2506,p2508,p2722,p2723);
FA fa84(p2717,p2510,p2514,p2724,p2725);
HA ha1278(p2719,p2721,p2726,p2727);
HA ha1279(p2516,p2518,p2728,p2729);
HA ha1280(p2520,p2723,p2730,p2731);
FA fa85(p2727,p2512,p2522,p2732,p2733);
FA fa86(p2524,p2526,p2725,p2734,p2735);
FA fa87(p2729,p2731,p2528,p2736,p2737);
FA fa88(p2530,p2532,p2534,p2738,p2739);
FA fa89(p2536,p2538,p2540,p2740,p2741);
HA ha1281(p2542,p2733,p2742,p2743);
FA fa90(p2735,p2737,p2544,p2744,p2745);
HA ha1282(p2546,p2548,p2746,p2747);
FA fa91(p2739,p2743,p2552,p2748,p2749);
HA ha1283(p2554,p2556,p2750,p2751);
HA ha1284(p2741,p2745,p2752,p2753);
FA fa92(p2747,p2550,p2558,p2754,p2755);
HA ha1285(p2560,p2562,p2756,p2757);
HA ha1286(p2749,p2751,p2758,p2759);
FA fa93(p2753,p2564,p2566,p2760,p2761);
FA fa94(p2568,p2570,p2757,p2762,p2763);
HA ha1287(p2759,p2574,p2764,p2765);
FA fa95(p2576,p2578,p2580,p2766,p2767);
FA fa96(p2755,p2582,p2584,p2768,p2769);
FA fa97(p2586,p2588,p2590,p2770,p2771);
HA ha1288(p2761,p2763,p2772,p2773);
HA ha1289(p2765,p2572,p2774,p2775);
HA ha1290(p2592,p2594,p2776,p2777);
FA fa98(p2596,p2598,p2767,p2778,p2779);
HA ha1291(p2773,p2602,p2780,p2781);
HA ha1292(p2604,p2769,p2782,p2783);
HA ha1293(p2771,p2775,p2784,p2785);
FA fa99(p2777,p2600,p2606,p2786,p2787);
HA ha1294(p2608,p2610,p2788,p2789);
FA fa100(p2612,p2779,p2781,p2790,p2791);
HA ha1295(p2783,p2785,p2792,p2793);
HA ha1296(p2614,p2616,p2794,p2795);
FA fa101(p2618,p2789,p2793,p2796,p2797);
FA fa102(p2624,p2787,p2791,p2798,p2799);
HA ha1297(p2795,p2620,p2800,p2801);
FA fa103(p2626,p2628,p2630,p2802,p2803);
FA fa104(p2797,p2622,p2632,p2804,p2805);
FA fa105(p2634,p2636,p2799,p2806,p2807);
FA fa106(p2801,p2638,p2640,p2808,p2809);
HA ha1298(p2642,p2803,p2810,p2811);
FA fa107(p2644,p2646,p2648,p2812,p2813);
HA ha1299(p2805,p2807,p2814,p2815);
HA ha1300(p2811,p2650,p2816,p2817);
FA fa108(p2652,p2654,p2656,p2818,p2819);
FA fa109(p2809,p2815,p2658,p2820,p2821);
HA ha1301(p2660,p2662,p2822,p2823);
FA fa110(p2664,p2813,p2817,p2824,p2825);
HA ha1302(p2666,p2670,p2826,p2827);
FA fa111(p2819,p2821,p2823,p2828,p2829);
FA fa112(p2672,p2674,p2676,p2830,p2831);
HA ha1303(p2825,p2827,p2832,p2833);
FA fa113(p2668,p2678,p2680,p2834,p2835);
HA ha1304(p2682,p2829,p2836,p2837);
FA fa114(p2833,p2684,p2686,p2838,p2839);
FA fa115(p2688,p2831,p2837,p2840,p2841);
HA ha1305(p2690,p2692,p2842,p2843);
HA ha1306(p2694,p2835,p2844,p2845);
FA fa116(p2696,p2698,p2839,p2846,p2847);
FA fa117(p2841,p2843,p2845,p2848,p2849);
FA fa118(p2700,p2702,p2704,p2850,p2851);
FA fa119(p2847,p2849,p2851,p2852,p2853);
HA ha1307(ip_11_15,ip_12_14,p2854,p2855);
FA fa120(ip_13_13,ip_14_12,ip_15_11,p2856,p2857);
FA fa121(p2706,p2708,p2710,p2858,p2859);
HA ha1308(p2855,p2712,p2860,p2861);
FA fa122(p2714,p2857,p2716,p2862,p2863);
FA fa123(p2859,p2861,p2720,p2864,p2865);
HA ha1309(p2863,p2718,p2866,p2867);
HA ha1310(p2726,p2865,p2868,p2869);
HA ha1311(p2722,p2728,p2870,p2871);
HA ha1312(p2730,p2867,p2872,p2873);
HA ha1313(p2869,p2724,p2874,p2875);
HA ha1314(p2871,p2873,p2876,p2877);
FA fa124(p2875,p2877,p2732,p2878,p2879);
FA fa125(p2734,p2736,p2742,p2880,p2881);
FA fa126(p2738,p2746,p2879,p2882,p2883);
FA fa127(p2740,p2744,p2750,p2884,p2885);
FA fa128(p2752,p2881,p2748,p2886,p2887);
HA ha1315(p2756,p2758,p2888,p2889);
FA fa129(p2883,p2885,p2887,p2890,p2891);
HA ha1316(p2889,p2754,p2892,p2893);
HA ha1317(p2764,p2760,p2894,p2895);
HA ha1318(p2762,p2772,p2896,p2897);
FA fa130(p2891,p2893,p2766,p2898,p2899);
FA fa131(p2774,p2776,p2895,p2900,p2901);
HA ha1319(p2897,p2768,p2902,p2903);
HA ha1320(p2770,p2780,p2904,p2905);
HA ha1321(p2782,p2784,p2906,p2907);
HA ha1322(p2899,p2778,p2908,p2909);
FA fa132(p2788,p2792,p2901,p2910,p2911);
HA ha1323(p2903,p2905,p2912,p2913);
FA fa133(p2907,p2794,p2909,p2914,p2915);
FA fa134(p2913,p2786,p2790,p2916,p2917);
HA ha1324(p2911,p2796,p2918,p2919);
FA fa135(p2800,p2915,p2798,p2920,p2921);
HA ha1325(p2917,p2919,p2922,p2923);
HA ha1326(p2802,p2810,p2924,p2925);
FA fa136(p2921,p2923,p2804,p2926,p2927);
FA fa137(p2806,p2814,p2925,p2928,p2929);
HA ha1327(p2808,p2816,p2930,p2931);
FA fa138(p2927,p2812,p2822,p2932,p2933);
FA fa139(p2929,p2931,p2818,p2934,p2935);
FA fa140(p2820,p2826,p2824,p2936,p2937);
HA ha1328(p2832,p2933,p2938,p2939);
FA fa141(p2935,p2828,p2836,p2940,p2941);
HA ha1329(p2937,p2939,p2942,p2943);
FA fa142(p2830,p2943,p2834,p2944,p2945);
FA fa143(p2842,p2844,p2941,p2946,p2947);
HA ha1330(p2838,p2840,p2948,p2949);
HA ha1331(p2945,p2947,p2950,p2951);
FA fa144(p2949,p2846,p2848,p2952,p2953);
HA ha1332(p2951,p2850,p2954,p2955);
HA ha1333(p2852,p2953,p2956,p2957);
FA fa145(ip_12_15,ip_13_14,ip_14_13,p2958,p2959);
HA ha1334(ip_15_12,p2854,p2960,p2961);
FA fa146(p2959,p2961,p2856,p2962,p2963);
HA ha1335(p2860,p2858,p2964,p2965);
FA fa147(p2963,p2862,p2965,p2966,p2967);
HA ha1336(p2864,p2866,p2968,p2969);
HA ha1337(p2868,p2870,p2970,p2971);
FA fa148(p2872,p2967,p2969,p2972,p2973);
HA ha1338(p2874,p2876,p2974,p2975);
HA ha1339(p2971,p2973,p2976,p2977);
FA fa149(p2975,p2977,p2878,p2978,p2979);
FA fa150(p2880,p2979,p2882,p2980,p2981);
FA fa151(p2888,p2884,p2886,p2982,p2983);
FA fa152(p2981,p2892,p2890,p2984,p2985);
FA fa153(p2894,p2896,p2983,p2986,p2987);
HA ha1340(p2985,p2898,p2988,p2989);
FA fa154(p2902,p2904,p2906,p2990,p2991);
HA ha1341(p2987,p2900,p2992,p2993);
HA ha1342(p2908,p2912,p2994,p2995);
FA fa155(p2989,p2991,p2993,p2996,p2997);
HA ha1343(p2995,p2910,p2998,p2999);
FA fa156(p2914,p2918,p2997,p3000,p3001);
FA fa157(p2999,p2916,p2922,p3002,p3003);
FA fa158(p2920,p2924,p3001,p3004,p3005);
FA fa159(p3003,p2926,p2930,p3006,p3007);
HA ha1344(p3005,p2928,p3008,p3009);
HA ha1345(p3007,p3009,p3010,p3011);
FA fa160(p2932,p2934,p2938,p3012,p3013);
HA ha1346(p3011,p2936,p3014,p3015);
FA fa161(p2942,p3013,p3015,p3016,p3017);
HA ha1347(p2940,p2944,p3018,p3019);
FA fa162(p2948,p3017,p2946,p3020,p3021);
FA fa163(p2950,p3019,p3021,p3022,p3023);
FA fa164(p2954,p3023,p2952,p3024,p3025);
HA ha1348(ip_13_15,ip_14_14,p3026,p3027);
HA ha1349(ip_15_13,p3027,p3028,p3029);
FA fa165(p2960,p3029,p2958,p3030,p3031);
FA fa166(p3031,p2962,p2964,p3032,p3033);
FA fa167(p2968,p3033,p2966,p3034,p3035);
FA fa168(p2970,p2974,p3035,p3036,p3037);
HA ha1350(p2972,p2976,p3038,p3039);
HA ha1351(p3037,p3039,p3040,p3041);
FA fa169(p3041,p2978,p2980,p3042,p3043);
HA ha1352(p3043,p2982,p3044,p3045);
HA ha1353(p2984,p3045,p3046,p3047);
FA fa170(p2986,p2988,p3047,p3048,p3049);
FA fa171(p2992,p2994,p2990,p3050,p3051);
FA fa172(p3049,p2998,p3051,p3052,p3053);
FA fa173(p2996,p3053,p3000,p3054,p3055);
FA fa174(p3002,p3055,p3004,p3056,p3057);
HA ha1354(p3008,p3057,p3058,p3059);
HA ha1355(p3006,p3010,p3060,p3061);
FA fa175(p3059,p3061,p3014,p3062,p3063);
HA ha1356(p3012,p3063,p3064,p3065);
HA ha1357(p3065,p3016,p3066,p3067);
HA ha1358(p3018,p3067,p3068,p3069);
FA fa176(p3020,p3069,p3022,p3070,p3071);
FA fa177(ip_14_15,ip_15_14,p3026,p3072,p3073);
FA fa178(p3028,p3073,p3030,p3074,p3075);
HA ha1359(p3075,p3032,p3076,p3077);
HA ha1360(p3077,p3034,p3078,p3079);
HA ha1361(p3038,p3079,p3080,p3081);
FA fa179(p3036,p3040,p3081,p3082,p3083);
FA fa180(p3083,p3042,p3044,p3084,p3085);
HA ha1362(p3046,p3085,p3086,p3087);
HA ha1363(p3087,p3048,p3088,p3089);
FA fa181(p3050,p3089,p3052,p3090,p3091);
FA fa182(p3091,p3054,p3056,p3092,p3093);
FA fa183(p3058,p3060,p3093,p3094,p3095);
HA ha1364(p3095,p3062,p3096,p3097);
FA fa184(p3064,p3097,p3066,p3098,p3099);
FA fa185(p3068,p3099,p3070,p3100,p3101);
FA fa186(ip_15_15,p3072,p3074,p3102,p3103);
FA fa187(p3103,p3076,p3078,p3104,p3105);
HA ha1365(p3080,p3105,p3106,p3107);
HA ha1366(p3107,p3082,p3108,p3109);
HA ha1367(p3109,p3084,p3110,p3111);
HA ha1368(p3086,p3111,p3112,p3113);
HA ha1369(p3113,p3088,p3114,p3115);
HA ha1370(p3115,p3090,p3116,p3117);
HA ha1371(p3117,p3092,p3118,p3119);
FA fa188(p3119,p3094,p3096,p3120,p3121);
FA fa189(p3121,p3098,p3100,p3122,p3123);
wire [31:0] a,b;
wire [31:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = ip_2_0;
assign b[2] = p1;
assign a[3] = p5;
assign b[3] = p7;
assign a[4] = p17;
assign b[4] = p19;
assign a[5] = p37;
assign b[5] = p39;
assign a[6] = p67;
assign b[6] = p69;
assign a[7] = p107;
assign b[7] = p105;
assign a[8] = p153;
assign b[8] = p155;
assign a[9] = p213;
assign b[9] = 1'b0;
assign a[10] = p212;
assign b[10] = p283;
assign a[11] = p367;
assign b[11] = p369;
assign a[12] = p463;
assign b[12] = p465;
assign a[13] = p577;
assign b[13] = 1'b0;
assign a[14] = p576;
assign b[14] = p707;
assign a[15] = p855;
assign b[15] = 1'b0;
assign a[16] = p1025;
assign b[16] = p854;
assign a[17] = p1205;
assign b[17] = p1207;
assign a[18] = p1403;
assign b[18] = p1405;
assign a[19] = p1609;
assign b[19] = p1611;
assign a[20] = p1823;
assign b[20] = p1825;
assign a[21] = p2043;
assign b[21] = p2045;
assign a[22] = p2269;
assign b[22] = p2271;
assign a[23] = p2489;
assign b[23] = p2491;
assign a[24] = p2703;
assign b[24] = p2705;
assign a[25] = p2853;
assign b[25] = 1'b0;
assign a[26] = p2955;
assign b[26] = p2957;
assign a[27] = p2956;
assign b[27] = p3025;
assign a[28] = p3071;
assign b[28] = p3024;
assign a[29] = p3101;
assign b[29] = 1'b0;
assign a[30] = p3123;
assign b[30] = 1'b0;
assign a[31] = p3102;
assign b[31] = p3104;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[31] = s[31] & p3106 & p3108 & p3110 & p3112 & p3114 & p3116 & p3118 & p3120 & p3122;
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 
// 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 
module adder(a,b,s);
input [31:0] a,b;
output [31:0] s;
wire c2,p0_0,g27_24,p1_1,g3_2,g27_26,g16_16,p27_26,g31_28,g21_20,g1_0,g24_24,g19_19,p30_30,g23_0,p23_22,p11_8,g29_28,p31_30,p25_24,c8,c11,g23_20,c25,g5_0,p6_6,c13,g15_8,g8_8,g19_0,p20_20,p8_8,p18_18,p9_9,p2_2,c9,c27,g20_20,g25_0,p7_7,p27_27,p31_16,p28_28,p24_24,p13_13,g31_30,g4_4,g31_16,c7,g11_8,c18,c21,g7_4,g28_28,c22,c26,c30,p10_10,g25_24,p15_14,p3_3,p7_6,c19,c0,g25_25,g0_0,c12,p23_20,g29_29,p12_12,g2_2,c14,p19_18,g27_27,g30_30,g17_16,g31_24,p25_25,p4_4,c5,g7_7,c4,c23,p9_8,g11_10,g13_12,p31_24,g10_10,p5_5,g23_16,g23_23,p7_4,g26_26,g29_0,g7_6,p17_17,g18_18,g11_0,g9_8,g15_14,g3_3,p17_16,c20,p31_31,c15,c29,g19_16,p11_10,g19_18,g17_17,g13_13,p27_24,g15_0,c16,g5_5,g21_21,p19_16,p29_29,g22_22,p14_14,g11_11,g9_0,g9_9,c17,g15_12,p5_4,g31_31,g12_12,c3,g17_0,g13_0,c1,g6_6,p29_28,c6,c24,p19_19,p11_11,p23_16,c28,p26_26,g5_4,p31_28,p15_12,g21_0,p22_22,p13_12,g27_0,p16_16,g23_22,p3_2,g14_14,p15_15,p23_23,g7_0,c31,p21_21,p21_20,g3_0,c10,g15_15,p15_8,g1_1;

assign p0_0 = a[0] ^ b[0];
assign g0_0 = a[0] & b[0];
assign p1_1 = a[1] ^ b[1];
assign g1_1 = a[1] & b[1];
assign p2_2 = a[2] ^ b[2];
assign g2_2 = a[2] & b[2];
assign p3_3 = a[3] ^ b[3];
assign g3_3 = a[3] & b[3];
assign p4_4 = a[4] ^ b[4];
assign g4_4 = a[4] & b[4];
assign p5_5 = a[5] ^ b[5];
assign g5_5 = a[5] & b[5];
assign p6_6 = a[6] ^ b[6];
assign g6_6 = a[6] & b[6];
assign p7_7 = a[7] ^ b[7];
assign g7_7 = a[7] & b[7];
assign p8_8 = a[8] ^ b[8];
assign g8_8 = a[8] & b[8];
assign p9_9 = a[9] ^ b[9];
assign g9_9 = a[9] & b[9];
assign p10_10 = a[10] ^ b[10];
assign g10_10 = a[10] & b[10];
assign p11_11 = a[11] ^ b[11];
assign g11_11 = a[11] & b[11];
assign p12_12 = a[12] ^ b[12];
assign g12_12 = a[12] & b[12];
assign p13_13 = a[13] ^ b[13];
assign g13_13 = a[13] & b[13];
assign p14_14 = a[14] ^ b[14];
assign g14_14 = a[14] & b[14];
assign p15_15 = a[15] ^ b[15];
assign g15_15 = a[15] & b[15];
assign p16_16 = a[16] ^ b[16];
assign g16_16 = a[16] & b[16];
assign p17_17 = a[17] ^ b[17];
assign g17_17 = a[17] & b[17];
assign p18_18 = a[18] ^ b[18];
assign g18_18 = a[18] & b[18];
assign p19_19 = a[19] ^ b[19];
assign g19_19 = a[19] & b[19];
assign p20_20 = a[20] ^ b[20];
assign g20_20 = a[20] & b[20];
assign p21_21 = a[21] ^ b[21];
assign g21_21 = a[21] & b[21];
assign p22_22 = a[22] ^ b[22];
assign g22_22 = a[22] & b[22];
assign p23_23 = a[23] ^ b[23];
assign g23_23 = a[23] & b[23];
assign p24_24 = a[24] ^ b[24];
assign g24_24 = a[24] & b[24];
assign p25_25 = a[25] ^ b[25];
assign g25_25 = a[25] & b[25];
assign p26_26 = a[26] ^ b[26];
assign g26_26 = a[26] & b[26];
assign p27_27 = a[27] ^ b[27];
assign g27_27 = a[27] & b[27];
assign p28_28 = a[28] ^ b[28];
assign g28_28 = a[28] & b[28];
assign p29_29 = a[29] ^ b[29];
assign g29_29 = a[29] & b[29];
assign p30_30 = a[30] ^ b[30];
assign g30_30 = a[30] & b[30];
assign p31_31 = a[31] ^ b[31];
assign g31_31 = a[31] & b[31];
assign g1_0 = c1;
assign g2_0 = c2;
assign g3_0 = c3;
assign g4_0 = c4;
assign g5_0 = c5;
assign g6_0 = c6;
assign g7_0 = c7;
assign g8_0 = c8;
assign g9_0 = c9;
assign g10_0 = c10;
assign g11_0 = c11;
assign g12_0 = c12;
assign g13_0 = c13;
assign g14_0 = c14;
assign g15_0 = c15;
assign g16_0 = c16;
assign g17_0 = c17;
assign g18_0 = c18;
assign g19_0 = c19;
assign g20_0 = c20;
assign g21_0 = c21;
assign g22_0 = c22;
assign g23_0 = c23;
assign g24_0 = c24;
assign g25_0 = c25;
assign g26_0 = c26;
assign g27_0 = c27;
assign g28_0 = c28;
assign g29_0 = c29;
assign g30_0 = c30;
assign g31_0 = c31;
BLACK black31_30(g31_31, p31_31, g30_30, p30_30, g31_30, p31_30);
BLACK black31_28(g31_30, p31_30, g29_28, p29_28, g31_28, p31_28);
BLACK black31_24(g31_28, p31_28, g27_24, p27_24, g31_24, p31_24);
BLACK black31_16(g31_24, p31_24, g23_16, p23_16, g31_16, p31_16);
GREY grey31(g31_16, p31_16, g15_0, c31);
GREY grey30(g30_30, p30_30, g29_0, c30);
BLACK black29_28(g29_29, p29_29, g28_28, p28_28, g29_28, p29_28);
GREY grey29(g29_28, p29_28, g27_0, c29);
GREY grey28(g28_28, p28_28, g27_0, c28);
BLACK black27_26(g27_27, p27_27, g26_26, p26_26, g27_26, p27_26);
BLACK black27_24(g27_26, p27_26, g25_24, p25_24, g27_24, p27_24);
GREY grey27(g27_24, p27_24, g23_0, c27);
GREY grey26(g26_26, p26_26, g25_0, c26);
BLACK black25_24(g25_25, p25_25, g24_24, p24_24, g25_24, p25_24);
GREY grey25(g25_24, p25_24, g23_0, c25);
GREY grey24(g24_24, p24_24, g23_0, c24);
BLACK black23_22(g23_23, p23_23, g22_22, p22_22, g23_22, p23_22);
BLACK black23_20(g23_22, p23_22, g21_20, p21_20, g23_20, p23_20);
BLACK black23_16(g23_20, p23_20, g19_16, p19_16, g23_16, p23_16);
GREY grey23(g23_16, p23_16, g15_0, c23);
GREY grey22(g22_22, p22_22, g21_0, c22);
BLACK black21_20(g21_21, p21_21, g20_20, p20_20, g21_20, p21_20);
GREY grey21(g21_20, p21_20, g19_0, c21);
GREY grey20(g20_20, p20_20, g19_0, c20);
BLACK black19_18(g19_19, p19_19, g18_18, p18_18, g19_18, p19_18);
BLACK black19_16(g19_18, p19_18, g17_16, p17_16, g19_16, p19_16);
GREY grey19(g19_16, p19_16, g15_0, c19);
GREY grey18(g18_18, p18_18, g17_0, c18);
BLACK black17_16(g17_17, p17_17, g16_16, p16_16, g17_16, p17_16);
GREY grey17(g17_16, p17_16, g15_0, c17);
GREY grey16(g16_16, p16_16, g15_0, c16);
BLACK black15_14(g15_15, p15_15, g14_14, p14_14, g15_14, p15_14);
BLACK black15_12(g15_14, p15_14, g13_12, p13_12, g15_12, p15_12);
BLACK black15_8(g15_12, p15_12, g11_8, p11_8, g15_8, p15_8);
GREY grey15(g15_8, p15_8, g7_0, c15);
GREY grey14(g14_14, p14_14, g13_0, c14);
BLACK black13_12(g13_13, p13_13, g12_12, p12_12, g13_12, p13_12);
GREY grey13(g13_12, p13_12, g11_0, c13);
GREY grey12(g12_12, p12_12, g11_0, c12);
BLACK black11_10(g11_11, p11_11, g10_10, p10_10, g11_10, p11_10);
BLACK black11_8(g11_10, p11_10, g9_8, p9_8, g11_8, p11_8);
GREY grey11(g11_8, p11_8, g7_0, c11);
GREY grey10(g10_10, p10_10, g9_0, c10);
BLACK black9_8(g9_9, p9_9, g8_8, p8_8, g9_8, p9_8);
GREY grey9(g9_8, p9_8, g7_0, c9);
GREY grey8(g8_8, p8_8, g7_0, c8);
BLACK black7_6(g7_7, p7_7, g6_6, p6_6, g7_6, p7_6);
BLACK black7_4(g7_6, p7_6, g5_4, p5_4, g7_4, p7_4);
GREY grey7(g7_4, p7_4, g3_0, c7);
GREY grey6(g6_6, p6_6, g5_0, c6);
BLACK black5_4(g5_5, p5_5, g4_4, p4_4, g5_4, p5_4);
GREY grey5(g5_4, p5_4, g3_0, c5);
GREY grey4(g4_4, p4_4, g3_0, c4);
BLACK black3_2(g3_3, p3_3, g2_2, p2_2, g3_2, p3_2);
GREY grey3(g3_2, p3_2, g1_0, c3);
GREY grey2(g2_2, p2_2, g1_0, c2);
GREY grey1(g1_1, p1_1, g0_0, c1);
assign s[0] = a[0] ^ b[0];
assign c0 = g0_0;
assign s[1] = p1_1 ^ c0;
assign s[2] = p2_2 ^ c1;
assign s[3] = p3_3 ^ c2;
assign s[4] = p4_4 ^ c3;
assign s[5] = p5_5 ^ c4;
assign s[6] = p6_6 ^ c5;
assign s[7] = p7_7 ^ c6;
assign s[8] = p8_8 ^ c7;
assign s[9] = p9_9 ^ c8;
assign s[10] = p10_10 ^ c9;
assign s[11] = p11_11 ^ c10;
assign s[12] = p12_12 ^ c11;
assign s[13] = p13_13 ^ c12;
assign s[14] = p14_14 ^ c13;
assign s[15] = p15_15 ^ c14;
assign s[16] = p16_16 ^ c15;
assign s[17] = p17_17 ^ c16;
assign s[18] = p18_18 ^ c17;
assign s[19] = p19_19 ^ c18;
assign s[20] = p20_20 ^ c19;
assign s[21] = p21_21 ^ c20;
assign s[22] = p22_22 ^ c21;
assign s[23] = p23_23 ^ c22;
assign s[24] = p24_24 ^ c23;
assign s[25] = p25_25 ^ c24;
assign s[26] = p26_26 ^ c25;
assign s[27] = p27_27 ^ c26;
assign s[28] = p28_28 ^ c27;
assign s[29] = p29_29 ^ c28;
assign s[30] = p30_30 ^ c29;
assign s[31] = p31_31 ^ c30;
endmodule

module GREY(gik, pik, gkj, gij);
input gik, pik, gkj;
output gij;
assign gij = gik | (pik & gkj);
endmodule

module BLACK(gik, pik, gkj, pkj, gij, pij);
input gik, pik, gkj, pkj;
output gij, pij;
assign pij = pik & pkj;
assign gij = gik | (pik & gkj);
endmodule

