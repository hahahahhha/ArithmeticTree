// 1 2 2 1 2 2 2 2 1 1 2 1 1 2 1 3 

module main(x,y,o);
input [7:0] x,y;
output [15:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_1_0,x[1],y[0]);
and and9(ip_1_1,x[1],y[1]);
and and10(ip_1_2,x[1],y[2]);
and and11(ip_1_3,x[1],y[3]);
and and12(ip_1_4,x[1],y[4]);
and and13(ip_1_5,x[1],y[5]);
and and14(ip_1_6,x[1],y[6]);
and and15(ip_1_7,x[1],y[7]);
and and16(ip_2_0,x[2],y[0]);
and and17(ip_2_1,x[2],y[1]);
and and18(ip_2_2,x[2],y[2]);
and and19(ip_2_3,x[2],y[3]);
and and20(ip_2_4,x[2],y[4]);
and and21(ip_2_5,x[2],y[5]);
and and22(ip_2_6,x[2],y[6]);
and and23(ip_2_7,x[2],y[7]);
and and24(ip_3_0,x[3],y[0]);
and and25(ip_3_1,x[3],y[1]);
and and26(ip_3_2,x[3],y[2]);
and and27(ip_3_3,x[3],y[3]);
and and28(ip_3_4,x[3],y[4]);
and and29(ip_3_5,x[3],y[5]);
and and30(ip_3_6,x[3],y[6]);
and and31(ip_3_7,x[3],y[7]);
and and32(ip_4_0,x[4],y[0]);
and and33(ip_4_1,x[4],y[1]);
and and34(ip_4_2,x[4],y[2]);
and and35(ip_4_3,x[4],y[3]);
and and36(ip_4_4,x[4],y[4]);
and and37(ip_4_5,x[4],y[5]);
and and38(ip_4_6,x[4],y[6]);
and and39(ip_4_7,x[4],y[7]);
and and40(ip_5_0,x[5],y[0]);
and and41(ip_5_1,x[5],y[1]);
and and42(ip_5_2,x[5],y[2]);
and and43(ip_5_3,x[5],y[3]);
and and44(ip_5_4,x[5],y[4]);
and and45(ip_5_5,x[5],y[5]);
and and46(ip_5_6,x[5],y[6]);
and and47(ip_5_7,x[5],y[7]);
and and48(ip_6_0,x[6],y[0]);
and and49(ip_6_1,x[6],y[1]);
and and50(ip_6_2,x[6],y[2]);
and and51(ip_6_3,x[6],y[3]);
and and52(ip_6_4,x[6],y[4]);
and and53(ip_6_5,x[6],y[5]);
and and54(ip_6_6,x[6],y[6]);
and and55(ip_6_7,x[6],y[7]);
and and56(ip_7_0,x[7],y[0]);
and and57(ip_7_1,x[7],y[1]);
and and58(ip_7_2,x[7],y[2]);
and and59(ip_7_3,x[7],y[3]);
and and60(ip_7_4,x[7],y[4]);
and and61(ip_7_5,x[7],y[5]);
and and62(ip_7_6,x[7],y[6]);
and and63(ip_7_7,x[7],y[7]);
HA ha0(ip_0_2,ip_1_1,p0,p1);
FA fa0(ip_0_3,ip_1_2,ip_2_1,p2,p3);
FA fa1(ip_3_0,p0,p3,p4,p5);
HA ha1(ip_0_4,ip_1_3,p6,p7);
FA fa2(ip_2_2,ip_3_1,ip_4_0,p8,p9);
HA ha2(p7,p9,p10,p11);
HA ha3(p11,p2,p12,p13);
FA fa3(ip_0_5,ip_1_4,ip_2_3,p14,p15);
FA fa4(ip_3_2,ip_4_1,ip_5_0,p16,p17);
HA ha4(p6,p15,p18,p19);
FA fa5(p17,p10,p19,p20,p21);
HA ha5(p8,p12,p22,p23);
FA fa6(ip_0_6,ip_1_5,ip_2_4,p24,p25);
HA ha6(ip_3_3,ip_4_2,p26,p27);
HA ha7(ip_5_1,ip_6_0,p28,p29);
HA ha8(p27,p29,p30,p31);
FA fa7(p25,p31,p14,p32,p33);
HA ha9(p16,p18,p34,p35);
FA fa8(p33,p35,p22,p36,p37);
FA fa9(ip_0_7,ip_1_6,ip_2_5,p38,p39);
FA fa10(ip_3_4,ip_4_3,ip_5_2,p40,p41);
FA fa11(ip_6_1,ip_7_0,p26,p42,p43);
FA fa12(p28,p30,p39,p44,p45);
FA fa13(p41,p43,p24,p46,p47);
HA ha10(p34,p45,p48,p49);
FA fa14(p47,p32,p49,p50,p51);
FA fa15(ip_1_7,ip_2_6,ip_3_5,p52,p53);
FA fa16(ip_4_4,ip_5_3,ip_6_2,p54,p55);
FA fa17(ip_7_1,p53,p55,p56,p57);
FA fa18(p38,p40,p42,p58,p59);
HA ha11(p57,p44,p60,p61);
HA ha12(p46,p48,p62,p63);
HA ha13(p59,p61,p64,p65);
FA fa19(p63,p65,p50,p66,p67);
HA ha14(ip_2_7,ip_3_6,p68,p69);
FA fa20(ip_4_5,ip_5_4,ip_6_3,p70,p71);
HA ha15(ip_7_2,p69,p72,p73);
HA ha16(p71,p73,p74,p75);
FA fa21(p52,p54,p75,p76,p77);
FA fa22(p56,p77,p58,p78,p79);
HA ha17(p60,p62,p80,p81);
HA ha18(p64,p79,p82,p83);
FA fa23(p81,p83,p66,p84,p85);
HA ha19(ip_3_7,ip_4_6,p86,p87);
HA ha20(ip_5_5,ip_6_4,p88,p89);
HA ha21(ip_7_3,p68,p90,p91);
FA fa24(p87,p89,p72,p92,p93);
FA fa25(p91,p70,p74,p94,p95);
HA ha22(p93,p95,p96,p97);
FA fa26(p76,p97,p80,p98,p99);
FA fa27(p78,p82,p99,p100,p101);
HA ha23(ip_4_7,ip_5_6,p102,p103);
FA fa28(ip_6_5,ip_7_4,p103,p104,p105);
FA fa29(p86,p88,p105,p106,p107);
HA ha24(p90,p107,p108,p109);
HA ha25(p109,p92,p110,p111);
HA ha26(p111,p94,p112,p113);
HA ha27(p96,p113,p114,p115);
FA fa30(p115,p98,p100,p116,p117);
HA ha28(ip_5_7,ip_6_6,p118,p119);
FA fa31(ip_7_5,p102,p119,p120,p121);
HA ha29(p104,p121,p122,p123);
HA ha30(p106,p108,p124,p125);
HA ha31(p123,p110,p126,p127);
HA ha32(p125,p127,p128,p129);
HA ha33(p112,p129,p130,p131);
FA fa32(p114,p131,p116,p132,p133);
HA ha34(ip_6_7,ip_7_6,p134,p135);
FA fa33(p118,p135,p120,p136,p137);
HA ha35(p122,p124,p138,p139);
FA fa34(p137,p126,p139,p140,p141);
FA fa35(p128,p130,p141,p142,p143);
HA ha36(ip_7_7,p134,p144,p145);
FA fa36(p145,p136,p138,p146,p147);
FA fa37(p147,p140,p142,p148,p149);
wire [15:0] a,b;
wire [15:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = ip_2_0;
assign b[2] = p1;
assign a[3] = p5;
assign b[3] = 1'b0;
assign a[4] = p13;
assign b[4] = p4;
assign a[5] = p21;
assign b[5] = p23;
assign a[6] = p20;
assign b[6] = p37;
assign a[7] = p36;
assign b[7] = p51;
assign a[8] = p67;
assign b[8] = 1'b0;
assign a[9] = p85;
assign b[9] = 1'b0;
assign a[10] = p101;
assign b[10] = p84;
assign a[11] = p117;
assign b[11] = 1'b0;
assign a[12] = p133;
assign b[12] = 1'b0;
assign a[13] = p143;
assign b[13] = p132;
assign a[14] = p149;
assign b[14] = 1'b0;
assign a[15] = p144;
assign b[15] = p146;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[15] = s[15] & p148;
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [15:0] a,b;
output [15:0] s;
assign s = a+b;
endmodule
