// 1 2 1 1 2 1 1 2 1 1 2 2 2 1 1 1 2 2 2 2 2 2 2 2 1 2 1 1 2 1 1 1 

module main(x,y,o);
input [15:0] x,y;
output [31:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_1_0,x[1],y[0]);
and and17(ip_1_1,x[1],y[1]);
and and18(ip_1_2,x[1],y[2]);
and and19(ip_1_3,x[1],y[3]);
and and20(ip_1_4,x[1],y[4]);
and and21(ip_1_5,x[1],y[5]);
and and22(ip_1_6,x[1],y[6]);
and and23(ip_1_7,x[1],y[7]);
and and24(ip_1_8,x[1],y[8]);
and and25(ip_1_9,x[1],y[9]);
and and26(ip_1_10,x[1],y[10]);
and and27(ip_1_11,x[1],y[11]);
and and28(ip_1_12,x[1],y[12]);
and and29(ip_1_13,x[1],y[13]);
and and30(ip_1_14,x[1],y[14]);
and and31(ip_1_15,x[1],y[15]);
and and32(ip_2_0,x[2],y[0]);
and and33(ip_2_1,x[2],y[1]);
and and34(ip_2_2,x[2],y[2]);
and and35(ip_2_3,x[2],y[3]);
and and36(ip_2_4,x[2],y[4]);
and and37(ip_2_5,x[2],y[5]);
and and38(ip_2_6,x[2],y[6]);
and and39(ip_2_7,x[2],y[7]);
and and40(ip_2_8,x[2],y[8]);
and and41(ip_2_9,x[2],y[9]);
and and42(ip_2_10,x[2],y[10]);
and and43(ip_2_11,x[2],y[11]);
and and44(ip_2_12,x[2],y[12]);
and and45(ip_2_13,x[2],y[13]);
and and46(ip_2_14,x[2],y[14]);
and and47(ip_2_15,x[2],y[15]);
and and48(ip_3_0,x[3],y[0]);
and and49(ip_3_1,x[3],y[1]);
and and50(ip_3_2,x[3],y[2]);
and and51(ip_3_3,x[3],y[3]);
and and52(ip_3_4,x[3],y[4]);
and and53(ip_3_5,x[3],y[5]);
and and54(ip_3_6,x[3],y[6]);
and and55(ip_3_7,x[3],y[7]);
and and56(ip_3_8,x[3],y[8]);
and and57(ip_3_9,x[3],y[9]);
and and58(ip_3_10,x[3],y[10]);
and and59(ip_3_11,x[3],y[11]);
and and60(ip_3_12,x[3],y[12]);
and and61(ip_3_13,x[3],y[13]);
and and62(ip_3_14,x[3],y[14]);
and and63(ip_3_15,x[3],y[15]);
and and64(ip_4_0,x[4],y[0]);
and and65(ip_4_1,x[4],y[1]);
and and66(ip_4_2,x[4],y[2]);
and and67(ip_4_3,x[4],y[3]);
and and68(ip_4_4,x[4],y[4]);
and and69(ip_4_5,x[4],y[5]);
and and70(ip_4_6,x[4],y[6]);
and and71(ip_4_7,x[4],y[7]);
and and72(ip_4_8,x[4],y[8]);
and and73(ip_4_9,x[4],y[9]);
and and74(ip_4_10,x[4],y[10]);
and and75(ip_4_11,x[4],y[11]);
and and76(ip_4_12,x[4],y[12]);
and and77(ip_4_13,x[4],y[13]);
and and78(ip_4_14,x[4],y[14]);
and and79(ip_4_15,x[4],y[15]);
and and80(ip_5_0,x[5],y[0]);
and and81(ip_5_1,x[5],y[1]);
and and82(ip_5_2,x[5],y[2]);
and and83(ip_5_3,x[5],y[3]);
and and84(ip_5_4,x[5],y[4]);
and and85(ip_5_5,x[5],y[5]);
and and86(ip_5_6,x[5],y[6]);
and and87(ip_5_7,x[5],y[7]);
and and88(ip_5_8,x[5],y[8]);
and and89(ip_5_9,x[5],y[9]);
and and90(ip_5_10,x[5],y[10]);
and and91(ip_5_11,x[5],y[11]);
and and92(ip_5_12,x[5],y[12]);
and and93(ip_5_13,x[5],y[13]);
and and94(ip_5_14,x[5],y[14]);
and and95(ip_5_15,x[5],y[15]);
and and96(ip_6_0,x[6],y[0]);
and and97(ip_6_1,x[6],y[1]);
and and98(ip_6_2,x[6],y[2]);
and and99(ip_6_3,x[6],y[3]);
and and100(ip_6_4,x[6],y[4]);
and and101(ip_6_5,x[6],y[5]);
and and102(ip_6_6,x[6],y[6]);
and and103(ip_6_7,x[6],y[7]);
and and104(ip_6_8,x[6],y[8]);
and and105(ip_6_9,x[6],y[9]);
and and106(ip_6_10,x[6],y[10]);
and and107(ip_6_11,x[6],y[11]);
and and108(ip_6_12,x[6],y[12]);
and and109(ip_6_13,x[6],y[13]);
and and110(ip_6_14,x[6],y[14]);
and and111(ip_6_15,x[6],y[15]);
and and112(ip_7_0,x[7],y[0]);
and and113(ip_7_1,x[7],y[1]);
and and114(ip_7_2,x[7],y[2]);
and and115(ip_7_3,x[7],y[3]);
and and116(ip_7_4,x[7],y[4]);
and and117(ip_7_5,x[7],y[5]);
and and118(ip_7_6,x[7],y[6]);
and and119(ip_7_7,x[7],y[7]);
and and120(ip_7_8,x[7],y[8]);
and and121(ip_7_9,x[7],y[9]);
and and122(ip_7_10,x[7],y[10]);
and and123(ip_7_11,x[7],y[11]);
and and124(ip_7_12,x[7],y[12]);
and and125(ip_7_13,x[7],y[13]);
and and126(ip_7_14,x[7],y[14]);
and and127(ip_7_15,x[7],y[15]);
and and128(ip_8_0,x[8],y[0]);
and and129(ip_8_1,x[8],y[1]);
and and130(ip_8_2,x[8],y[2]);
and and131(ip_8_3,x[8],y[3]);
and and132(ip_8_4,x[8],y[4]);
and and133(ip_8_5,x[8],y[5]);
and and134(ip_8_6,x[8],y[6]);
and and135(ip_8_7,x[8],y[7]);
and and136(ip_8_8,x[8],y[8]);
and and137(ip_8_9,x[8],y[9]);
and and138(ip_8_10,x[8],y[10]);
and and139(ip_8_11,x[8],y[11]);
and and140(ip_8_12,x[8],y[12]);
and and141(ip_8_13,x[8],y[13]);
and and142(ip_8_14,x[8],y[14]);
and and143(ip_8_15,x[8],y[15]);
and and144(ip_9_0,x[9],y[0]);
and and145(ip_9_1,x[9],y[1]);
and and146(ip_9_2,x[9],y[2]);
and and147(ip_9_3,x[9],y[3]);
and and148(ip_9_4,x[9],y[4]);
and and149(ip_9_5,x[9],y[5]);
and and150(ip_9_6,x[9],y[6]);
and and151(ip_9_7,x[9],y[7]);
and and152(ip_9_8,x[9],y[8]);
and and153(ip_9_9,x[9],y[9]);
and and154(ip_9_10,x[9],y[10]);
and and155(ip_9_11,x[9],y[11]);
and and156(ip_9_12,x[9],y[12]);
and and157(ip_9_13,x[9],y[13]);
and and158(ip_9_14,x[9],y[14]);
and and159(ip_9_15,x[9],y[15]);
and and160(ip_10_0,x[10],y[0]);
and and161(ip_10_1,x[10],y[1]);
and and162(ip_10_2,x[10],y[2]);
and and163(ip_10_3,x[10],y[3]);
and and164(ip_10_4,x[10],y[4]);
and and165(ip_10_5,x[10],y[5]);
and and166(ip_10_6,x[10],y[6]);
and and167(ip_10_7,x[10],y[7]);
and and168(ip_10_8,x[10],y[8]);
and and169(ip_10_9,x[10],y[9]);
and and170(ip_10_10,x[10],y[10]);
and and171(ip_10_11,x[10],y[11]);
and and172(ip_10_12,x[10],y[12]);
and and173(ip_10_13,x[10],y[13]);
and and174(ip_10_14,x[10],y[14]);
and and175(ip_10_15,x[10],y[15]);
and and176(ip_11_0,x[11],y[0]);
and and177(ip_11_1,x[11],y[1]);
and and178(ip_11_2,x[11],y[2]);
and and179(ip_11_3,x[11],y[3]);
and and180(ip_11_4,x[11],y[4]);
and and181(ip_11_5,x[11],y[5]);
and and182(ip_11_6,x[11],y[6]);
and and183(ip_11_7,x[11],y[7]);
and and184(ip_11_8,x[11],y[8]);
and and185(ip_11_9,x[11],y[9]);
and and186(ip_11_10,x[11],y[10]);
and and187(ip_11_11,x[11],y[11]);
and and188(ip_11_12,x[11],y[12]);
and and189(ip_11_13,x[11],y[13]);
and and190(ip_11_14,x[11],y[14]);
and and191(ip_11_15,x[11],y[15]);
and and192(ip_12_0,x[12],y[0]);
and and193(ip_12_1,x[12],y[1]);
and and194(ip_12_2,x[12],y[2]);
and and195(ip_12_3,x[12],y[3]);
and and196(ip_12_4,x[12],y[4]);
and and197(ip_12_5,x[12],y[5]);
and and198(ip_12_6,x[12],y[6]);
and and199(ip_12_7,x[12],y[7]);
and and200(ip_12_8,x[12],y[8]);
and and201(ip_12_9,x[12],y[9]);
and and202(ip_12_10,x[12],y[10]);
and and203(ip_12_11,x[12],y[11]);
and and204(ip_12_12,x[12],y[12]);
and and205(ip_12_13,x[12],y[13]);
and and206(ip_12_14,x[12],y[14]);
and and207(ip_12_15,x[12],y[15]);
and and208(ip_13_0,x[13],y[0]);
and and209(ip_13_1,x[13],y[1]);
and and210(ip_13_2,x[13],y[2]);
and and211(ip_13_3,x[13],y[3]);
and and212(ip_13_4,x[13],y[4]);
and and213(ip_13_5,x[13],y[5]);
and and214(ip_13_6,x[13],y[6]);
and and215(ip_13_7,x[13],y[7]);
and and216(ip_13_8,x[13],y[8]);
and and217(ip_13_9,x[13],y[9]);
and and218(ip_13_10,x[13],y[10]);
and and219(ip_13_11,x[13],y[11]);
and and220(ip_13_12,x[13],y[12]);
and and221(ip_13_13,x[13],y[13]);
and and222(ip_13_14,x[13],y[14]);
and and223(ip_13_15,x[13],y[15]);
and and224(ip_14_0,x[14],y[0]);
and and225(ip_14_1,x[14],y[1]);
and and226(ip_14_2,x[14],y[2]);
and and227(ip_14_3,x[14],y[3]);
and and228(ip_14_4,x[14],y[4]);
and and229(ip_14_5,x[14],y[5]);
and and230(ip_14_6,x[14],y[6]);
and and231(ip_14_7,x[14],y[7]);
and and232(ip_14_8,x[14],y[8]);
and and233(ip_14_9,x[14],y[9]);
and and234(ip_14_10,x[14],y[10]);
and and235(ip_14_11,x[14],y[11]);
and and236(ip_14_12,x[14],y[12]);
and and237(ip_14_13,x[14],y[13]);
and and238(ip_14_14,x[14],y[14]);
and and239(ip_14_15,x[14],y[15]);
and and240(ip_15_0,x[15],y[0]);
and and241(ip_15_1,x[15],y[1]);
and and242(ip_15_2,x[15],y[2]);
and and243(ip_15_3,x[15],y[3]);
and and244(ip_15_4,x[15],y[4]);
and and245(ip_15_5,x[15],y[5]);
and and246(ip_15_6,x[15],y[6]);
and and247(ip_15_7,x[15],y[7]);
and and248(ip_15_8,x[15],y[8]);
and and249(ip_15_9,x[15],y[9]);
and and250(ip_15_10,x[15],y[10]);
and and251(ip_15_11,x[15],y[11]);
and and252(ip_15_12,x[15],y[12]);
and and253(ip_15_13,x[15],y[13]);
and and254(ip_15_14,x[15],y[14]);
and and255(ip_15_15,x[15],y[15]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
FA fa2(ip_3_0,p3,p0,p4,p5);
FA fa3(ip_0_4,ip_1_3,ip_2_2,p6,p7);
HA ha0(ip_3_1,ip_4_0,p8,p9);
FA fa4(p9,p7,p2,p10,p11);
FA fa5(ip_0_5,ip_1_4,ip_2_3,p12,p13);
FA fa6(ip_3_2,ip_4_1,ip_5_0,p14,p15);
FA fa7(p8,p13,p15,p16,p17);
FA fa8(p6,p17,p10,p18,p19);
FA fa9(ip_0_6,ip_1_5,ip_2_4,p20,p21);
FA fa10(ip_3_3,ip_4_2,ip_5_1,p22,p23);
FA fa11(ip_6_0,p21,p23,p24,p25);
FA fa12(p12,p14,p25,p26,p27);
FA fa13(p16,p27,p18,p28,p29);
FA fa14(ip_0_7,ip_1_6,ip_2_5,p30,p31);
HA ha1(ip_3_4,ip_4_3,p32,p33);
FA fa15(ip_5_2,ip_6_1,ip_7_0,p34,p35);
FA fa16(p33,p31,p35,p36,p37);
FA fa17(p20,p22,p37,p38,p39);
FA fa18(p24,p39,p26,p40,p41);
FA fa19(ip_0_8,ip_1_7,ip_2_6,p42,p43);
HA ha2(ip_3_5,ip_4_4,p44,p45);
FA fa20(ip_5_3,ip_6_2,ip_7_1,p46,p47);
HA ha3(ip_8_0,p32,p48,p49);
FA fa21(p45,p43,p47,p50,p51);
FA fa22(p49,p30,p34,p52,p53);
FA fa23(p51,p36,p53,p54,p55);
FA fa24(p38,p55,p40,p56,p57);
FA fa25(ip_0_9,ip_1_8,ip_2_7,p58,p59);
FA fa26(ip_3_6,ip_4_5,ip_5_4,p60,p61);
HA ha4(ip_6_3,ip_7_2,p62,p63);
FA fa27(ip_8_1,ip_9_0,p44,p64,p65);
FA fa28(p63,p48,p59,p66,p67);
FA fa29(p61,p65,p42,p68,p69);
FA fa30(p46,p67,p69,p70,p71);
FA fa31(p50,p52,p71,p72,p73);
FA fa32(p54,p73,p56,p74,p75);
FA fa33(ip_0_10,ip_1_9,ip_2_8,p76,p77);
FA fa34(ip_3_7,ip_4_6,ip_5_5,p78,p79);
HA ha5(ip_6_4,ip_7_3,p80,p81);
FA fa35(ip_8_2,ip_9_1,ip_10_0,p82,p83);
FA fa36(p62,p81,p77,p84,p85);
HA ha6(p79,p83,p86,p87);
FA fa37(p58,p60,p64,p88,p89);
FA fa38(p85,p87,p66,p90,p91);
FA fa39(p68,p89,p91,p92,p93);
FA fa40(p70,p93,p72,p94,p95);
FA fa41(ip_0_11,ip_1_10,ip_2_9,p96,p97);
FA fa42(ip_3_8,ip_4_7,ip_5_6,p98,p99);
FA fa43(ip_6_5,ip_7_4,ip_8_3,p100,p101);
FA fa44(ip_9_2,ip_10_1,ip_11_0,p102,p103);
FA fa45(p80,p101,p103,p104,p105);
FA fa46(p97,p99,p76,p106,p107);
FA fa47(p78,p82,p86,p108,p109);
FA fa48(p105,p107,p84,p110,p111);
FA fa49(p109,p111,p88,p112,p113);
FA fa50(p90,p113,p92,p114,p115);
FA fa51(ip_0_12,ip_1_11,ip_2_10,p116,p117);
FA fa52(ip_3_9,ip_4_8,ip_5_7,p118,p119);
FA fa53(ip_6_6,ip_7_5,ip_8_4,p120,p121);
FA fa54(ip_9_3,ip_10_2,ip_11_1,p122,p123);
FA fa55(ip_12_0,p117,p119,p124,p125);
HA ha7(p121,p123,p126,p127);
FA fa56(p100,p102,p127,p128,p129);
FA fa57(p96,p98,p125,p130,p131);
FA fa58(p104,p106,p129,p132,p133);
FA fa59(p131,p108,p110,p134,p135);
FA fa60(p133,p135,p112,p136,p137);
FA fa61(ip_0_13,ip_1_12,ip_2_11,p138,p139);
FA fa62(ip_3_10,ip_4_9,ip_5_8,p140,p141);
FA fa63(ip_6_7,ip_7_6,ip_8_5,p142,p143);
FA fa64(ip_9_4,ip_10_3,ip_11_2,p144,p145);
FA fa65(ip_12_1,ip_13_0,p139,p146,p147);
FA fa66(p141,p143,p145,p148,p149);
FA fa67(p116,p118,p120,p150,p151);
FA fa68(p122,p126,p147,p152,p153);
FA fa69(p149,p124,p151,p154,p155);
FA fa70(p153,p128,p130,p156,p157);
FA fa71(p155,p132,p157,p158,p159);
FA fa72(p134,p159,p136,p160,p161);
FA fa73(ip_0_14,ip_1_13,ip_2_12,p162,p163);
FA fa74(ip_3_11,ip_4_10,ip_5_9,p164,p165);
FA fa75(ip_6_8,ip_7_7,ip_8_6,p166,p167);
FA fa76(ip_9_5,ip_10_4,ip_11_3,p168,p169);
FA fa77(ip_12_2,ip_13_1,ip_14_0,p170,p171);
FA fa78(p163,p165,p167,p172,p173);
FA fa79(p169,p171,p138,p174,p175);
FA fa80(p140,p142,p144,p176,p177);
FA fa81(p146,p173,p175,p178,p179);
FA fa82(p148,p177,p150,p180,p181);
FA fa83(p152,p179,p181,p182,p183);
FA fa84(p154,p183,p156,p184,p185);
FA fa85(p185,p158,p160,p186,p187);
FA fa86(ip_0_15,ip_1_14,ip_2_13,p188,p189);
FA fa87(ip_3_12,ip_4_11,ip_5_10,p190,p191);
HA ha8(ip_6_9,ip_7_8,p192,p193);
FA fa88(ip_8_7,ip_9_6,ip_10_5,p194,p195);
FA fa89(ip_11_4,ip_12_3,ip_13_2,p196,p197);
FA fa90(ip_14_1,ip_15_0,p193,p198,p199);
FA fa91(p189,p191,p195,p200,p201);
FA fa92(p197,p199,p162,p202,p203);
FA fa93(p164,p166,p168,p204,p205);
FA fa94(p170,p201,p203,p206,p207);
HA ha9(p172,p174,p208,p209);
FA fa95(p205,p176,p207,p210,p211);
FA fa96(p209,p178,p180,p212,p213);
FA fa97(p211,p182,p213,p214,p215);
FA fa98(p184,p215,p186,p216,p217);
HA ha10(ip_1_15,ip_2_14,p218,p219);
FA fa99(ip_3_13,ip_4_12,ip_5_11,p220,p221);
FA fa100(ip_6_10,ip_7_9,ip_8_8,p222,p223);
FA fa101(ip_9_7,ip_10_6,ip_11_5,p224,p225);
FA fa102(ip_12_4,ip_13_3,ip_14_2,p226,p227);
FA fa103(ip_15_1,p192,p219,p228,p229);
FA fa104(p221,p223,p225,p230,p231);
FA fa105(p227,p188,p190,p232,p233);
FA fa106(p194,p196,p198,p234,p235);
FA fa107(p229,p231,p200,p236,p237);
HA ha11(p202,p233,p238,p239);
FA fa108(p235,p204,p208,p240,p241);
FA fa109(p237,p239,p206,p242,p243);
FA fa110(p241,p243,p210,p244,p245);
FA fa111(p212,p245,p214,p246,p247);
FA fa112(ip_2_15,ip_3_14,ip_4_13,p248,p249);
FA fa113(ip_5_12,ip_6_11,ip_7_10,p250,p251);
FA fa114(ip_8_9,ip_9_8,ip_10_7,p252,p253);
FA fa115(ip_11_6,ip_12_5,ip_13_4,p254,p255);
FA fa116(ip_14_3,ip_15_2,p218,p256,p257);
FA fa117(p249,p251,p253,p258,p259);
FA fa118(p255,p257,p220,p260,p261);
FA fa119(p222,p224,p226,p262,p263);
FA fa120(p228,p259,p261,p264,p265);
FA fa121(p230,p263,p232,p266,p267);
FA fa122(p234,p238,p265,p268,p269);
FA fa123(p236,p267,p269,p270,p271);
FA fa124(p240,p242,p271,p272,p273);
HA ha12(p244,p273,p274,p275);
FA fa125(ip_3_15,ip_4_14,ip_5_13,p276,p277);
FA fa126(ip_6_12,ip_7_11,ip_8_10,p278,p279);
FA fa127(ip_9_9,ip_10_8,ip_11_7,p280,p281);
FA fa128(ip_12_6,ip_13_5,ip_14_4,p282,p283);
FA fa129(ip_15_3,p277,p279,p284,p285);
FA fa130(p281,p283,p248,p286,p287);
HA ha13(p250,p252,p288,p289);
FA fa131(p254,p256,p285,p290,p291);
FA fa132(p287,p289,p258,p292,p293);
FA fa133(p260,p291,p262,p294,p295);
FA fa134(p293,p264,p295,p296,p297);
FA fa135(p266,p268,p297,p298,p299);
HA ha14(p270,p299,p300,p301);
HA ha15(p272,p274,p302,p303);
FA fa136(ip_4_15,ip_5_14,ip_6_13,p304,p305);
FA fa137(ip_7_12,ip_8_11,ip_9_10,p306,p307);
FA fa138(ip_10_9,ip_11_8,ip_12_7,p308,p309);
FA fa139(ip_13_6,ip_14_5,ip_15_4,p310,p311);
FA fa140(p305,p307,p309,p312,p313);
FA fa141(p311,p276,p278,p314,p315);
FA fa142(p280,p282,p288,p316,p317);
FA fa143(p313,p284,p286,p318,p319);
FA fa144(p315,p317,p290,p320,p321);
FA fa145(p292,p319,p321,p322,p323);
FA fa146(p294,p323,p296,p324,p325);
FA fa147(p325,p298,p300,p326,p327);
FA fa148(ip_5_15,ip_6_14,ip_7_13,p328,p329);
FA fa149(ip_8_12,ip_9_11,ip_10_10,p330,p331);
FA fa150(ip_11_9,ip_12_8,ip_13_7,p332,p333);
FA fa151(ip_14_6,ip_15_5,p329,p334,p335);
FA fa152(p331,p333,p304,p336,p337);
HA ha16(p306,p308,p338,p339);
FA fa153(p310,p335,p337,p340,p341);
HA ha17(p339,p312,p342,p343);
HA ha18(p341,p314,p344,p345);
FA fa154(p316,p343,p345,p346,p347);
FA fa155(p318,p320,p347,p348,p349);
FA fa156(p322,p349,p324,p350,p351);
FA fa157(ip_6_15,ip_7_14,ip_8_13,p352,p353);
FA fa158(ip_9_12,ip_10_11,ip_11_10,p354,p355);
FA fa159(ip_12_9,ip_13_8,ip_14_7,p356,p357);
FA fa160(ip_15_6,p353,p355,p358,p359);
HA ha19(p357,p328,p360,p361);
FA fa161(p330,p332,p334,p362,p363);
FA fa162(p338,p359,p361,p364,p365);
FA fa163(p336,p363,p340,p366,p367);
FA fa164(p342,p365,p344,p368,p369);
HA ha20(p367,p369,p370,p371);
FA fa165(p346,p371,p348,p372,p373);
FA fa166(ip_7_15,ip_8_14,ip_9_13,p374,p375);
FA fa167(ip_10_12,ip_11_11,ip_12_10,p376,p377);
FA fa168(ip_13_9,ip_14_8,ip_15_7,p378,p379);
FA fa169(p375,p377,p379,p380,p381);
FA fa170(p352,p354,p356,p382,p383);
FA fa171(p360,p381,p358,p384,p385);
FA fa172(p383,p362,p385,p386,p387);
FA fa173(p364,p366,p387,p388,p389);
FA fa174(p368,p370,p389,p390,p391);
FA fa175(ip_8_15,ip_9_14,ip_10_13,p392,p393);
FA fa176(ip_11_12,ip_12_11,ip_13_10,p394,p395);
HA ha21(ip_14_9,ip_15_8,p396,p397);
FA fa177(p397,p393,p395,p398,p399);
FA fa178(p374,p376,p378,p400,p401);
FA fa179(p399,p380,p401,p402,p403);
FA fa180(p382,p384,p403,p404,p405);
FA fa181(p386,p405,p388,p406,p407);
HA ha22(ip_9_15,ip_10_14,p408,p409);
HA ha23(ip_11_13,ip_12_12,p410,p411);
FA fa182(ip_13_11,ip_14_10,ip_15_9,p412,p413);
FA fa183(p396,p409,p411,p414,p415);
FA fa184(p413,p392,p394,p416,p417);
FA fa185(p415,p398,p417,p418,p419);
FA fa186(p400,p419,p402,p420,p421);
FA fa187(p421,p404,p406,p422,p423);
FA fa188(ip_10_15,ip_11_14,ip_12_13,p424,p425);
FA fa189(ip_13_12,ip_14_11,ip_15_10,p426,p427);
FA fa190(p408,p410,p425,p428,p429);
FA fa191(p427,p412,p429,p430,p431);
FA fa192(p414,p431,p416,p432,p433);
FA fa193(p433,p418,p420,p434,p435);
FA fa194(ip_11_15,ip_12_14,ip_13_13,p436,p437);
FA fa195(ip_14_12,ip_15_11,p437,p438,p439);
FA fa196(p424,p426,p439,p440,p441);
FA fa197(p428,p441,p430,p442,p443);
FA fa198(p443,p432,p434,p444,p445);
FA fa199(ip_12_15,ip_13_14,ip_14_13,p446,p447);
FA fa200(ip_15_12,p447,p436,p448,p449);
FA fa201(p438,p449,p440,p450,p451);
FA fa202(p451,p442,p444,p452,p453);
FA fa203(ip_13_15,ip_14_14,ip_15_13,p454,p455);
FA fa204(p455,p446,p448,p456,p457);
HA ha24(p457,p450,p458,p459);
FA fa205(ip_14_15,ip_15_14,p454,p460,p461);
FA fa206(p461,p456,p458,p462,p463);
FA fa207(ip_15_15,p460,p462,p464,p465);
wire [31:0] a,b;
wire [31:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p5;
assign b[3] = 1'b0;
assign a[4] = p11;
assign b[4] = p4;
assign a[5] = p19;
assign b[5] = 1'b0;
assign a[6] = p29;
assign b[6] = 1'b0;
assign a[7] = p41;
assign b[7] = p28;
assign a[8] = p57;
assign b[8] = 1'b0;
assign a[9] = p75;
assign b[9] = 1'b0;
assign a[10] = p95;
assign b[10] = p74;
assign a[11] = p115;
assign b[11] = p94;
assign a[12] = p137;
assign b[12] = p114;
assign a[13] = p161;
assign b[13] = 1'b0;
assign a[14] = p187;
assign b[14] = 1'b0;
assign a[15] = p217;
assign b[15] = 1'b0;
assign a[16] = p247;
assign b[16] = p216;
assign a[17] = p275;
assign b[17] = p246;
assign a[18] = p301;
assign b[18] = p303;
assign a[19] = p302;
assign b[19] = p327;
assign a[20] = p351;
assign b[20] = p326;
assign a[21] = p373;
assign b[21] = p350;
assign a[22] = p391;
assign b[22] = p372;
assign a[23] = p390;
assign b[23] = p407;
assign a[24] = p423;
assign b[24] = 1'b0;
assign a[25] = p435;
assign b[25] = p422;
assign a[26] = p445;
assign b[26] = 1'b0;
assign a[27] = p453;
assign b[27] = 1'b0;
assign a[28] = p459;
assign b[28] = p452;
assign a[29] = p463;
assign b[29] = 1'b0;
assign a[30] = p465;
assign b[30] = 1'b0;
assign a[31] = p464;
assign b[31] = 1'b0;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[31] = s[31];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [31:0] a,b;
output [31:0] s;
assign s = a+b;
endmodule
