// 1 2 1 1 1 1 1 2 1 1 2 2 2 2 2 2 1 1 2 1 1 2 1 1 2 1 2 2 1 1 2 2 2 1 2 2 1 1 1 2 2 1 1 2 2 1 2 1 1 2 1 1 2 2 2 2 1 1 2 2 1 1 2 1 

module main(x,y,o);
input [31:0] x,y;
output [63:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_0_16,ip_0_17,ip_0_18,ip_0_19,ip_0_20,ip_0_21,ip_0_22,ip_0_23,ip_0_24,ip_0_25,ip_0_26,ip_0_27,ip_0_28,ip_0_29,ip_0_30,ip_0_31,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_1_16,ip_1_17,ip_1_18,ip_1_19,ip_1_20,ip_1_21,ip_1_22,ip_1_23,ip_1_24,ip_1_25,ip_1_26,ip_1_27,ip_1_28,ip_1_29,ip_1_30,ip_1_31,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_2_16,ip_2_17,ip_2_18,ip_2_19,ip_2_20,ip_2_21,ip_2_22,ip_2_23,ip_2_24,ip_2_25,ip_2_26,ip_2_27,ip_2_28,ip_2_29,ip_2_30,ip_2_31,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_3_16,ip_3_17,ip_3_18,ip_3_19,ip_3_20,ip_3_21,ip_3_22,ip_3_23,ip_3_24,ip_3_25,ip_3_26,ip_3_27,ip_3_28,ip_3_29,ip_3_30,ip_3_31,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_4_16,ip_4_17,ip_4_18,ip_4_19,ip_4_20,ip_4_21,ip_4_22,ip_4_23,ip_4_24,ip_4_25,ip_4_26,ip_4_27,ip_4_28,ip_4_29,ip_4_30,ip_4_31,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_5_16,ip_5_17,ip_5_18,ip_5_19,ip_5_20,ip_5_21,ip_5_22,ip_5_23,ip_5_24,ip_5_25,ip_5_26,ip_5_27,ip_5_28,ip_5_29,ip_5_30,ip_5_31,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_6_16,ip_6_17,ip_6_18,ip_6_19,ip_6_20,ip_6_21,ip_6_22,ip_6_23,ip_6_24,ip_6_25,ip_6_26,ip_6_27,ip_6_28,ip_6_29,ip_6_30,ip_6_31,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_7_16,ip_7_17,ip_7_18,ip_7_19,ip_7_20,ip_7_21,ip_7_22,ip_7_23,ip_7_24,ip_7_25,ip_7_26,ip_7_27,ip_7_28,ip_7_29,ip_7_30,ip_7_31,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_8_16,ip_8_17,ip_8_18,ip_8_19,ip_8_20,ip_8_21,ip_8_22,ip_8_23,ip_8_24,ip_8_25,ip_8_26,ip_8_27,ip_8_28,ip_8_29,ip_8_30,ip_8_31,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_9_16,ip_9_17,ip_9_18,ip_9_19,ip_9_20,ip_9_21,ip_9_22,ip_9_23,ip_9_24,ip_9_25,ip_9_26,ip_9_27,ip_9_28,ip_9_29,ip_9_30,ip_9_31,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_10_16,ip_10_17,ip_10_18,ip_10_19,ip_10_20,ip_10_21,ip_10_22,ip_10_23,ip_10_24,ip_10_25,ip_10_26,ip_10_27,ip_10_28,ip_10_29,ip_10_30,ip_10_31,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_11_16,ip_11_17,ip_11_18,ip_11_19,ip_11_20,ip_11_21,ip_11_22,ip_11_23,ip_11_24,ip_11_25,ip_11_26,ip_11_27,ip_11_28,ip_11_29,ip_11_30,ip_11_31,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_12_16,ip_12_17,ip_12_18,ip_12_19,ip_12_20,ip_12_21,ip_12_22,ip_12_23,ip_12_24,ip_12_25,ip_12_26,ip_12_27,ip_12_28,ip_12_29,ip_12_30,ip_12_31,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_13_16,ip_13_17,ip_13_18,ip_13_19,ip_13_20,ip_13_21,ip_13_22,ip_13_23,ip_13_24,ip_13_25,ip_13_26,ip_13_27,ip_13_28,ip_13_29,ip_13_30,ip_13_31,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_14_16,ip_14_17,ip_14_18,ip_14_19,ip_14_20,ip_14_21,ip_14_22,ip_14_23,ip_14_24,ip_14_25,ip_14_26,ip_14_27,ip_14_28,ip_14_29,ip_14_30,ip_14_31,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15,ip_15_16,ip_15_17,ip_15_18,ip_15_19,ip_15_20,ip_15_21,ip_15_22,ip_15_23,ip_15_24,ip_15_25,ip_15_26,ip_15_27,ip_15_28,ip_15_29,ip_15_30,ip_15_31,ip_16_0,ip_16_1,ip_16_2,ip_16_3,ip_16_4,ip_16_5,ip_16_6,ip_16_7,ip_16_8,ip_16_9,ip_16_10,ip_16_11,ip_16_12,ip_16_13,ip_16_14,ip_16_15,ip_16_16,ip_16_17,ip_16_18,ip_16_19,ip_16_20,ip_16_21,ip_16_22,ip_16_23,ip_16_24,ip_16_25,ip_16_26,ip_16_27,ip_16_28,ip_16_29,ip_16_30,ip_16_31,ip_17_0,ip_17_1,ip_17_2,ip_17_3,ip_17_4,ip_17_5,ip_17_6,ip_17_7,ip_17_8,ip_17_9,ip_17_10,ip_17_11,ip_17_12,ip_17_13,ip_17_14,ip_17_15,ip_17_16,ip_17_17,ip_17_18,ip_17_19,ip_17_20,ip_17_21,ip_17_22,ip_17_23,ip_17_24,ip_17_25,ip_17_26,ip_17_27,ip_17_28,ip_17_29,ip_17_30,ip_17_31,ip_18_0,ip_18_1,ip_18_2,ip_18_3,ip_18_4,ip_18_5,ip_18_6,ip_18_7,ip_18_8,ip_18_9,ip_18_10,ip_18_11,ip_18_12,ip_18_13,ip_18_14,ip_18_15,ip_18_16,ip_18_17,ip_18_18,ip_18_19,ip_18_20,ip_18_21,ip_18_22,ip_18_23,ip_18_24,ip_18_25,ip_18_26,ip_18_27,ip_18_28,ip_18_29,ip_18_30,ip_18_31,ip_19_0,ip_19_1,ip_19_2,ip_19_3,ip_19_4,ip_19_5,ip_19_6,ip_19_7,ip_19_8,ip_19_9,ip_19_10,ip_19_11,ip_19_12,ip_19_13,ip_19_14,ip_19_15,ip_19_16,ip_19_17,ip_19_18,ip_19_19,ip_19_20,ip_19_21,ip_19_22,ip_19_23,ip_19_24,ip_19_25,ip_19_26,ip_19_27,ip_19_28,ip_19_29,ip_19_30,ip_19_31,ip_20_0,ip_20_1,ip_20_2,ip_20_3,ip_20_4,ip_20_5,ip_20_6,ip_20_7,ip_20_8,ip_20_9,ip_20_10,ip_20_11,ip_20_12,ip_20_13,ip_20_14,ip_20_15,ip_20_16,ip_20_17,ip_20_18,ip_20_19,ip_20_20,ip_20_21,ip_20_22,ip_20_23,ip_20_24,ip_20_25,ip_20_26,ip_20_27,ip_20_28,ip_20_29,ip_20_30,ip_20_31,ip_21_0,ip_21_1,ip_21_2,ip_21_3,ip_21_4,ip_21_5,ip_21_6,ip_21_7,ip_21_8,ip_21_9,ip_21_10,ip_21_11,ip_21_12,ip_21_13,ip_21_14,ip_21_15,ip_21_16,ip_21_17,ip_21_18,ip_21_19,ip_21_20,ip_21_21,ip_21_22,ip_21_23,ip_21_24,ip_21_25,ip_21_26,ip_21_27,ip_21_28,ip_21_29,ip_21_30,ip_21_31,ip_22_0,ip_22_1,ip_22_2,ip_22_3,ip_22_4,ip_22_5,ip_22_6,ip_22_7,ip_22_8,ip_22_9,ip_22_10,ip_22_11,ip_22_12,ip_22_13,ip_22_14,ip_22_15,ip_22_16,ip_22_17,ip_22_18,ip_22_19,ip_22_20,ip_22_21,ip_22_22,ip_22_23,ip_22_24,ip_22_25,ip_22_26,ip_22_27,ip_22_28,ip_22_29,ip_22_30,ip_22_31,ip_23_0,ip_23_1,ip_23_2,ip_23_3,ip_23_4,ip_23_5,ip_23_6,ip_23_7,ip_23_8,ip_23_9,ip_23_10,ip_23_11,ip_23_12,ip_23_13,ip_23_14,ip_23_15,ip_23_16,ip_23_17,ip_23_18,ip_23_19,ip_23_20,ip_23_21,ip_23_22,ip_23_23,ip_23_24,ip_23_25,ip_23_26,ip_23_27,ip_23_28,ip_23_29,ip_23_30,ip_23_31,ip_24_0,ip_24_1,ip_24_2,ip_24_3,ip_24_4,ip_24_5,ip_24_6,ip_24_7,ip_24_8,ip_24_9,ip_24_10,ip_24_11,ip_24_12,ip_24_13,ip_24_14,ip_24_15,ip_24_16,ip_24_17,ip_24_18,ip_24_19,ip_24_20,ip_24_21,ip_24_22,ip_24_23,ip_24_24,ip_24_25,ip_24_26,ip_24_27,ip_24_28,ip_24_29,ip_24_30,ip_24_31,ip_25_0,ip_25_1,ip_25_2,ip_25_3,ip_25_4,ip_25_5,ip_25_6,ip_25_7,ip_25_8,ip_25_9,ip_25_10,ip_25_11,ip_25_12,ip_25_13,ip_25_14,ip_25_15,ip_25_16,ip_25_17,ip_25_18,ip_25_19,ip_25_20,ip_25_21,ip_25_22,ip_25_23,ip_25_24,ip_25_25,ip_25_26,ip_25_27,ip_25_28,ip_25_29,ip_25_30,ip_25_31,ip_26_0,ip_26_1,ip_26_2,ip_26_3,ip_26_4,ip_26_5,ip_26_6,ip_26_7,ip_26_8,ip_26_9,ip_26_10,ip_26_11,ip_26_12,ip_26_13,ip_26_14,ip_26_15,ip_26_16,ip_26_17,ip_26_18,ip_26_19,ip_26_20,ip_26_21,ip_26_22,ip_26_23,ip_26_24,ip_26_25,ip_26_26,ip_26_27,ip_26_28,ip_26_29,ip_26_30,ip_26_31,ip_27_0,ip_27_1,ip_27_2,ip_27_3,ip_27_4,ip_27_5,ip_27_6,ip_27_7,ip_27_8,ip_27_9,ip_27_10,ip_27_11,ip_27_12,ip_27_13,ip_27_14,ip_27_15,ip_27_16,ip_27_17,ip_27_18,ip_27_19,ip_27_20,ip_27_21,ip_27_22,ip_27_23,ip_27_24,ip_27_25,ip_27_26,ip_27_27,ip_27_28,ip_27_29,ip_27_30,ip_27_31,ip_28_0,ip_28_1,ip_28_2,ip_28_3,ip_28_4,ip_28_5,ip_28_6,ip_28_7,ip_28_8,ip_28_9,ip_28_10,ip_28_11,ip_28_12,ip_28_13,ip_28_14,ip_28_15,ip_28_16,ip_28_17,ip_28_18,ip_28_19,ip_28_20,ip_28_21,ip_28_22,ip_28_23,ip_28_24,ip_28_25,ip_28_26,ip_28_27,ip_28_28,ip_28_29,ip_28_30,ip_28_31,ip_29_0,ip_29_1,ip_29_2,ip_29_3,ip_29_4,ip_29_5,ip_29_6,ip_29_7,ip_29_8,ip_29_9,ip_29_10,ip_29_11,ip_29_12,ip_29_13,ip_29_14,ip_29_15,ip_29_16,ip_29_17,ip_29_18,ip_29_19,ip_29_20,ip_29_21,ip_29_22,ip_29_23,ip_29_24,ip_29_25,ip_29_26,ip_29_27,ip_29_28,ip_29_29,ip_29_30,ip_29_31,ip_30_0,ip_30_1,ip_30_2,ip_30_3,ip_30_4,ip_30_5,ip_30_6,ip_30_7,ip_30_8,ip_30_9,ip_30_10,ip_30_11,ip_30_12,ip_30_13,ip_30_14,ip_30_15,ip_30_16,ip_30_17,ip_30_18,ip_30_19,ip_30_20,ip_30_21,ip_30_22,ip_30_23,ip_30_24,ip_30_25,ip_30_26,ip_30_27,ip_30_28,ip_30_29,ip_30_30,ip_30_31,ip_31_0,ip_31_1,ip_31_2,ip_31_3,ip_31_4,ip_31_5,ip_31_6,ip_31_7,ip_31_8,ip_31_9,ip_31_10,ip_31_11,ip_31_12,ip_31_13,ip_31_14,ip_31_15,ip_31_16,ip_31_17,ip_31_18,ip_31_19,ip_31_20,ip_31_21,ip_31_22,ip_31_23,ip_31_24,ip_31_25,ip_31_26,ip_31_27,ip_31_28,ip_31_29,ip_31_30,ip_31_31;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149,p1150,p1151,p1152,p1153,p1154,p1155,p1156,p1157,p1158,p1159,p1160,p1161,p1162,p1163,p1164,p1165,p1166,p1167,p1168,p1169,p1170,p1171,p1172,p1173,p1174,p1175,p1176,p1177,p1178,p1179,p1180,p1181,p1182,p1183,p1184,p1185,p1186,p1187,p1188,p1189,p1190,p1191,p1192,p1193,p1194,p1195,p1196,p1197,p1198,p1199,p1200,p1201,p1202,p1203,p1204,p1205,p1206,p1207,p1208,p1209,p1210,p1211,p1212,p1213,p1214,p1215,p1216,p1217,p1218,p1219,p1220,p1221,p1222,p1223,p1224,p1225,p1226,p1227,p1228,p1229,p1230,p1231,p1232,p1233,p1234,p1235,p1236,p1237,p1238,p1239,p1240,p1241,p1242,p1243,p1244,p1245,p1246,p1247,p1248,p1249,p1250,p1251,p1252,p1253,p1254,p1255,p1256,p1257,p1258,p1259,p1260,p1261,p1262,p1263,p1264,p1265,p1266,p1267,p1268,p1269,p1270,p1271,p1272,p1273,p1274,p1275,p1276,p1277,p1278,p1279,p1280,p1281,p1282,p1283,p1284,p1285,p1286,p1287,p1288,p1289,p1290,p1291,p1292,p1293,p1294,p1295,p1296,p1297,p1298,p1299,p1300,p1301,p1302,p1303,p1304,p1305,p1306,p1307,p1308,p1309,p1310,p1311,p1312,p1313,p1314,p1315,p1316,p1317,p1318,p1319,p1320,p1321,p1322,p1323,p1324,p1325,p1326,p1327,p1328,p1329,p1330,p1331,p1332,p1333,p1334,p1335,p1336,p1337,p1338,p1339,p1340,p1341,p1342,p1343,p1344,p1345,p1346,p1347,p1348,p1349,p1350,p1351,p1352,p1353,p1354,p1355,p1356,p1357,p1358,p1359,p1360,p1361,p1362,p1363,p1364,p1365,p1366,p1367,p1368,p1369,p1370,p1371,p1372,p1373,p1374,p1375,p1376,p1377,p1378,p1379,p1380,p1381,p1382,p1383,p1384,p1385,p1386,p1387,p1388,p1389,p1390,p1391,p1392,p1393,p1394,p1395,p1396,p1397,p1398,p1399,p1400,p1401,p1402,p1403,p1404,p1405,p1406,p1407,p1408,p1409,p1410,p1411,p1412,p1413,p1414,p1415,p1416,p1417,p1418,p1419,p1420,p1421,p1422,p1423,p1424,p1425,p1426,p1427,p1428,p1429,p1430,p1431,p1432,p1433,p1434,p1435,p1436,p1437,p1438,p1439,p1440,p1441,p1442,p1443,p1444,p1445,p1446,p1447,p1448,p1449,p1450,p1451,p1452,p1453,p1454,p1455,p1456,p1457,p1458,p1459,p1460,p1461,p1462,p1463,p1464,p1465,p1466,p1467,p1468,p1469,p1470,p1471,p1472,p1473,p1474,p1475,p1476,p1477,p1478,p1479,p1480,p1481,p1482,p1483,p1484,p1485,p1486,p1487,p1488,p1489,p1490,p1491,p1492,p1493,p1494,p1495,p1496,p1497,p1498,p1499,p1500,p1501,p1502,p1503,p1504,p1505,p1506,p1507,p1508,p1509,p1510,p1511,p1512,p1513,p1514,p1515,p1516,p1517,p1518,p1519,p1520,p1521,p1522,p1523,p1524,p1525,p1526,p1527,p1528,p1529,p1530,p1531,p1532,p1533,p1534,p1535,p1536,p1537,p1538,p1539,p1540,p1541,p1542,p1543,p1544,p1545,p1546,p1547,p1548,p1549,p1550,p1551,p1552,p1553,p1554,p1555,p1556,p1557,p1558,p1559,p1560,p1561,p1562,p1563,p1564,p1565,p1566,p1567,p1568,p1569,p1570,p1571,p1572,p1573,p1574,p1575,p1576,p1577,p1578,p1579,p1580,p1581,p1582,p1583,p1584,p1585,p1586,p1587,p1588,p1589,p1590,p1591,p1592,p1593,p1594,p1595,p1596,p1597,p1598,p1599,p1600,p1601,p1602,p1603,p1604,p1605,p1606,p1607,p1608,p1609,p1610,p1611,p1612,p1613,p1614,p1615,p1616,p1617,p1618,p1619,p1620,p1621,p1622,p1623,p1624,p1625,p1626,p1627,p1628,p1629,p1630,p1631,p1632,p1633,p1634,p1635,p1636,p1637,p1638,p1639,p1640,p1641,p1642,p1643,p1644,p1645,p1646,p1647,p1648,p1649,p1650,p1651,p1652,p1653,p1654,p1655,p1656,p1657,p1658,p1659,p1660,p1661,p1662,p1663,p1664,p1665,p1666,p1667,p1668,p1669,p1670,p1671,p1672,p1673,p1674,p1675,p1676,p1677,p1678,p1679,p1680,p1681,p1682,p1683,p1684,p1685,p1686,p1687,p1688,p1689,p1690,p1691,p1692,p1693,p1694,p1695,p1696,p1697,p1698,p1699,p1700,p1701,p1702,p1703,p1704,p1705,p1706,p1707,p1708,p1709,p1710,p1711,p1712,p1713,p1714,p1715,p1716,p1717,p1718,p1719,p1720,p1721,p1722,p1723,p1724,p1725,p1726,p1727,p1728,p1729,p1730,p1731,p1732,p1733,p1734,p1735,p1736,p1737,p1738,p1739,p1740,p1741,p1742,p1743,p1744,p1745,p1746,p1747,p1748,p1749,p1750,p1751,p1752,p1753,p1754,p1755,p1756,p1757,p1758,p1759,p1760,p1761,p1762,p1763,p1764,p1765,p1766,p1767,p1768,p1769,p1770,p1771,p1772,p1773,p1774,p1775,p1776,p1777,p1778,p1779,p1780,p1781,p1782,p1783,p1784,p1785,p1786,p1787,p1788,p1789,p1790,p1791,p1792,p1793,p1794,p1795,p1796,p1797,p1798,p1799,p1800,p1801,p1802,p1803,p1804,p1805,p1806,p1807,p1808,p1809,p1810,p1811,p1812,p1813,p1814,p1815,p1816,p1817,p1818,p1819,p1820,p1821,p1822,p1823,p1824,p1825,p1826,p1827,p1828,p1829,p1830,p1831,p1832,p1833,p1834,p1835,p1836,p1837,p1838,p1839,p1840,p1841,p1842,p1843,p1844,p1845,p1846,p1847,p1848,p1849,p1850,p1851,p1852,p1853,p1854,p1855,p1856,p1857,p1858,p1859,p1860,p1861,p1862,p1863,p1864,p1865,p1866,p1867,p1868,p1869,p1870,p1871,p1872,p1873,p1874,p1875,p1876,p1877,p1878,p1879,p1880,p1881,p1882,p1883,p1884,p1885,p1886,p1887,p1888,p1889,p1890,p1891,p1892,p1893,p1894,p1895,p1896,p1897,p1898,p1899,p1900,p1901,p1902,p1903,p1904,p1905,p1906,p1907,p1908,p1909,p1910,p1911,p1912,p1913,p1914,p1915,p1916,p1917,p1918,p1919,p1920,p1921,p1922,p1923,p1924,p1925,p1926,p1927,p1928,p1929,p1930,p1931,p1932,p1933,p1934,p1935,p1936,p1937,p1938,p1939,p1940,p1941,p1942,p1943,p1944,p1945,p1946,p1947,p1948,p1949,p1950,p1951,p1952,p1953,p1954,p1955,p1956,p1957,p1958,p1959,p1960,p1961,p1962,p1963,p1964,p1965,p1966,p1967,p1968,p1969,p1970,p1971,p1972,p1973,p1974,p1975,p1976,p1977,p1978,p1979,p1980,p1981,p1982,p1983,p1984,p1985,p1986,p1987,p1988,p1989,p1990,p1991,p1992,p1993,p1994,p1995,p1996,p1997,p1998,p1999,p2000,p2001,p2002,p2003,p2004,p2005,p2006,p2007;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_0_16,x[0],y[16]);
and and17(ip_0_17,x[0],y[17]);
and and18(ip_0_18,x[0],y[18]);
and and19(ip_0_19,x[0],y[19]);
and and20(ip_0_20,x[0],y[20]);
and and21(ip_0_21,x[0],y[21]);
and and22(ip_0_22,x[0],y[22]);
and and23(ip_0_23,x[0],y[23]);
and and24(ip_0_24,x[0],y[24]);
and and25(ip_0_25,x[0],y[25]);
and and26(ip_0_26,x[0],y[26]);
and and27(ip_0_27,x[0],y[27]);
and and28(ip_0_28,x[0],y[28]);
and and29(ip_0_29,x[0],y[29]);
and and30(ip_0_30,x[0],y[30]);
and and31(ip_0_31,x[0],y[31]);
and and32(ip_1_0,x[1],y[0]);
and and33(ip_1_1,x[1],y[1]);
and and34(ip_1_2,x[1],y[2]);
and and35(ip_1_3,x[1],y[3]);
and and36(ip_1_4,x[1],y[4]);
and and37(ip_1_5,x[1],y[5]);
and and38(ip_1_6,x[1],y[6]);
and and39(ip_1_7,x[1],y[7]);
and and40(ip_1_8,x[1],y[8]);
and and41(ip_1_9,x[1],y[9]);
and and42(ip_1_10,x[1],y[10]);
and and43(ip_1_11,x[1],y[11]);
and and44(ip_1_12,x[1],y[12]);
and and45(ip_1_13,x[1],y[13]);
and and46(ip_1_14,x[1],y[14]);
and and47(ip_1_15,x[1],y[15]);
and and48(ip_1_16,x[1],y[16]);
and and49(ip_1_17,x[1],y[17]);
and and50(ip_1_18,x[1],y[18]);
and and51(ip_1_19,x[1],y[19]);
and and52(ip_1_20,x[1],y[20]);
and and53(ip_1_21,x[1],y[21]);
and and54(ip_1_22,x[1],y[22]);
and and55(ip_1_23,x[1],y[23]);
and and56(ip_1_24,x[1],y[24]);
and and57(ip_1_25,x[1],y[25]);
and and58(ip_1_26,x[1],y[26]);
and and59(ip_1_27,x[1],y[27]);
and and60(ip_1_28,x[1],y[28]);
and and61(ip_1_29,x[1],y[29]);
and and62(ip_1_30,x[1],y[30]);
and and63(ip_1_31,x[1],y[31]);
and and64(ip_2_0,x[2],y[0]);
and and65(ip_2_1,x[2],y[1]);
and and66(ip_2_2,x[2],y[2]);
and and67(ip_2_3,x[2],y[3]);
and and68(ip_2_4,x[2],y[4]);
and and69(ip_2_5,x[2],y[5]);
and and70(ip_2_6,x[2],y[6]);
and and71(ip_2_7,x[2],y[7]);
and and72(ip_2_8,x[2],y[8]);
and and73(ip_2_9,x[2],y[9]);
and and74(ip_2_10,x[2],y[10]);
and and75(ip_2_11,x[2],y[11]);
and and76(ip_2_12,x[2],y[12]);
and and77(ip_2_13,x[2],y[13]);
and and78(ip_2_14,x[2],y[14]);
and and79(ip_2_15,x[2],y[15]);
and and80(ip_2_16,x[2],y[16]);
and and81(ip_2_17,x[2],y[17]);
and and82(ip_2_18,x[2],y[18]);
and and83(ip_2_19,x[2],y[19]);
and and84(ip_2_20,x[2],y[20]);
and and85(ip_2_21,x[2],y[21]);
and and86(ip_2_22,x[2],y[22]);
and and87(ip_2_23,x[2],y[23]);
and and88(ip_2_24,x[2],y[24]);
and and89(ip_2_25,x[2],y[25]);
and and90(ip_2_26,x[2],y[26]);
and and91(ip_2_27,x[2],y[27]);
and and92(ip_2_28,x[2],y[28]);
and and93(ip_2_29,x[2],y[29]);
and and94(ip_2_30,x[2],y[30]);
and and95(ip_2_31,x[2],y[31]);
and and96(ip_3_0,x[3],y[0]);
and and97(ip_3_1,x[3],y[1]);
and and98(ip_3_2,x[3],y[2]);
and and99(ip_3_3,x[3],y[3]);
and and100(ip_3_4,x[3],y[4]);
and and101(ip_3_5,x[3],y[5]);
and and102(ip_3_6,x[3],y[6]);
and and103(ip_3_7,x[3],y[7]);
and and104(ip_3_8,x[3],y[8]);
and and105(ip_3_9,x[3],y[9]);
and and106(ip_3_10,x[3],y[10]);
and and107(ip_3_11,x[3],y[11]);
and and108(ip_3_12,x[3],y[12]);
and and109(ip_3_13,x[3],y[13]);
and and110(ip_3_14,x[3],y[14]);
and and111(ip_3_15,x[3],y[15]);
and and112(ip_3_16,x[3],y[16]);
and and113(ip_3_17,x[3],y[17]);
and and114(ip_3_18,x[3],y[18]);
and and115(ip_3_19,x[3],y[19]);
and and116(ip_3_20,x[3],y[20]);
and and117(ip_3_21,x[3],y[21]);
and and118(ip_3_22,x[3],y[22]);
and and119(ip_3_23,x[3],y[23]);
and and120(ip_3_24,x[3],y[24]);
and and121(ip_3_25,x[3],y[25]);
and and122(ip_3_26,x[3],y[26]);
and and123(ip_3_27,x[3],y[27]);
and and124(ip_3_28,x[3],y[28]);
and and125(ip_3_29,x[3],y[29]);
and and126(ip_3_30,x[3],y[30]);
and and127(ip_3_31,x[3],y[31]);
and and128(ip_4_0,x[4],y[0]);
and and129(ip_4_1,x[4],y[1]);
and and130(ip_4_2,x[4],y[2]);
and and131(ip_4_3,x[4],y[3]);
and and132(ip_4_4,x[4],y[4]);
and and133(ip_4_5,x[4],y[5]);
and and134(ip_4_6,x[4],y[6]);
and and135(ip_4_7,x[4],y[7]);
and and136(ip_4_8,x[4],y[8]);
and and137(ip_4_9,x[4],y[9]);
and and138(ip_4_10,x[4],y[10]);
and and139(ip_4_11,x[4],y[11]);
and and140(ip_4_12,x[4],y[12]);
and and141(ip_4_13,x[4],y[13]);
and and142(ip_4_14,x[4],y[14]);
and and143(ip_4_15,x[4],y[15]);
and and144(ip_4_16,x[4],y[16]);
and and145(ip_4_17,x[4],y[17]);
and and146(ip_4_18,x[4],y[18]);
and and147(ip_4_19,x[4],y[19]);
and and148(ip_4_20,x[4],y[20]);
and and149(ip_4_21,x[4],y[21]);
and and150(ip_4_22,x[4],y[22]);
and and151(ip_4_23,x[4],y[23]);
and and152(ip_4_24,x[4],y[24]);
and and153(ip_4_25,x[4],y[25]);
and and154(ip_4_26,x[4],y[26]);
and and155(ip_4_27,x[4],y[27]);
and and156(ip_4_28,x[4],y[28]);
and and157(ip_4_29,x[4],y[29]);
and and158(ip_4_30,x[4],y[30]);
and and159(ip_4_31,x[4],y[31]);
and and160(ip_5_0,x[5],y[0]);
and and161(ip_5_1,x[5],y[1]);
and and162(ip_5_2,x[5],y[2]);
and and163(ip_5_3,x[5],y[3]);
and and164(ip_5_4,x[5],y[4]);
and and165(ip_5_5,x[5],y[5]);
and and166(ip_5_6,x[5],y[6]);
and and167(ip_5_7,x[5],y[7]);
and and168(ip_5_8,x[5],y[8]);
and and169(ip_5_9,x[5],y[9]);
and and170(ip_5_10,x[5],y[10]);
and and171(ip_5_11,x[5],y[11]);
and and172(ip_5_12,x[5],y[12]);
and and173(ip_5_13,x[5],y[13]);
and and174(ip_5_14,x[5],y[14]);
and and175(ip_5_15,x[5],y[15]);
and and176(ip_5_16,x[5],y[16]);
and and177(ip_5_17,x[5],y[17]);
and and178(ip_5_18,x[5],y[18]);
and and179(ip_5_19,x[5],y[19]);
and and180(ip_5_20,x[5],y[20]);
and and181(ip_5_21,x[5],y[21]);
and and182(ip_5_22,x[5],y[22]);
and and183(ip_5_23,x[5],y[23]);
and and184(ip_5_24,x[5],y[24]);
and and185(ip_5_25,x[5],y[25]);
and and186(ip_5_26,x[5],y[26]);
and and187(ip_5_27,x[5],y[27]);
and and188(ip_5_28,x[5],y[28]);
and and189(ip_5_29,x[5],y[29]);
and and190(ip_5_30,x[5],y[30]);
and and191(ip_5_31,x[5],y[31]);
and and192(ip_6_0,x[6],y[0]);
and and193(ip_6_1,x[6],y[1]);
and and194(ip_6_2,x[6],y[2]);
and and195(ip_6_3,x[6],y[3]);
and and196(ip_6_4,x[6],y[4]);
and and197(ip_6_5,x[6],y[5]);
and and198(ip_6_6,x[6],y[6]);
and and199(ip_6_7,x[6],y[7]);
and and200(ip_6_8,x[6],y[8]);
and and201(ip_6_9,x[6],y[9]);
and and202(ip_6_10,x[6],y[10]);
and and203(ip_6_11,x[6],y[11]);
and and204(ip_6_12,x[6],y[12]);
and and205(ip_6_13,x[6],y[13]);
and and206(ip_6_14,x[6],y[14]);
and and207(ip_6_15,x[6],y[15]);
and and208(ip_6_16,x[6],y[16]);
and and209(ip_6_17,x[6],y[17]);
and and210(ip_6_18,x[6],y[18]);
and and211(ip_6_19,x[6],y[19]);
and and212(ip_6_20,x[6],y[20]);
and and213(ip_6_21,x[6],y[21]);
and and214(ip_6_22,x[6],y[22]);
and and215(ip_6_23,x[6],y[23]);
and and216(ip_6_24,x[6],y[24]);
and and217(ip_6_25,x[6],y[25]);
and and218(ip_6_26,x[6],y[26]);
and and219(ip_6_27,x[6],y[27]);
and and220(ip_6_28,x[6],y[28]);
and and221(ip_6_29,x[6],y[29]);
and and222(ip_6_30,x[6],y[30]);
and and223(ip_6_31,x[6],y[31]);
and and224(ip_7_0,x[7],y[0]);
and and225(ip_7_1,x[7],y[1]);
and and226(ip_7_2,x[7],y[2]);
and and227(ip_7_3,x[7],y[3]);
and and228(ip_7_4,x[7],y[4]);
and and229(ip_7_5,x[7],y[5]);
and and230(ip_7_6,x[7],y[6]);
and and231(ip_7_7,x[7],y[7]);
and and232(ip_7_8,x[7],y[8]);
and and233(ip_7_9,x[7],y[9]);
and and234(ip_7_10,x[7],y[10]);
and and235(ip_7_11,x[7],y[11]);
and and236(ip_7_12,x[7],y[12]);
and and237(ip_7_13,x[7],y[13]);
and and238(ip_7_14,x[7],y[14]);
and and239(ip_7_15,x[7],y[15]);
and and240(ip_7_16,x[7],y[16]);
and and241(ip_7_17,x[7],y[17]);
and and242(ip_7_18,x[7],y[18]);
and and243(ip_7_19,x[7],y[19]);
and and244(ip_7_20,x[7],y[20]);
and and245(ip_7_21,x[7],y[21]);
and and246(ip_7_22,x[7],y[22]);
and and247(ip_7_23,x[7],y[23]);
and and248(ip_7_24,x[7],y[24]);
and and249(ip_7_25,x[7],y[25]);
and and250(ip_7_26,x[7],y[26]);
and and251(ip_7_27,x[7],y[27]);
and and252(ip_7_28,x[7],y[28]);
and and253(ip_7_29,x[7],y[29]);
and and254(ip_7_30,x[7],y[30]);
and and255(ip_7_31,x[7],y[31]);
and and256(ip_8_0,x[8],y[0]);
and and257(ip_8_1,x[8],y[1]);
and and258(ip_8_2,x[8],y[2]);
and and259(ip_8_3,x[8],y[3]);
and and260(ip_8_4,x[8],y[4]);
and and261(ip_8_5,x[8],y[5]);
and and262(ip_8_6,x[8],y[6]);
and and263(ip_8_7,x[8],y[7]);
and and264(ip_8_8,x[8],y[8]);
and and265(ip_8_9,x[8],y[9]);
and and266(ip_8_10,x[8],y[10]);
and and267(ip_8_11,x[8],y[11]);
and and268(ip_8_12,x[8],y[12]);
and and269(ip_8_13,x[8],y[13]);
and and270(ip_8_14,x[8],y[14]);
and and271(ip_8_15,x[8],y[15]);
and and272(ip_8_16,x[8],y[16]);
and and273(ip_8_17,x[8],y[17]);
and and274(ip_8_18,x[8],y[18]);
and and275(ip_8_19,x[8],y[19]);
and and276(ip_8_20,x[8],y[20]);
and and277(ip_8_21,x[8],y[21]);
and and278(ip_8_22,x[8],y[22]);
and and279(ip_8_23,x[8],y[23]);
and and280(ip_8_24,x[8],y[24]);
and and281(ip_8_25,x[8],y[25]);
and and282(ip_8_26,x[8],y[26]);
and and283(ip_8_27,x[8],y[27]);
and and284(ip_8_28,x[8],y[28]);
and and285(ip_8_29,x[8],y[29]);
and and286(ip_8_30,x[8],y[30]);
and and287(ip_8_31,x[8],y[31]);
and and288(ip_9_0,x[9],y[0]);
and and289(ip_9_1,x[9],y[1]);
and and290(ip_9_2,x[9],y[2]);
and and291(ip_9_3,x[9],y[3]);
and and292(ip_9_4,x[9],y[4]);
and and293(ip_9_5,x[9],y[5]);
and and294(ip_9_6,x[9],y[6]);
and and295(ip_9_7,x[9],y[7]);
and and296(ip_9_8,x[9],y[8]);
and and297(ip_9_9,x[9],y[9]);
and and298(ip_9_10,x[9],y[10]);
and and299(ip_9_11,x[9],y[11]);
and and300(ip_9_12,x[9],y[12]);
and and301(ip_9_13,x[9],y[13]);
and and302(ip_9_14,x[9],y[14]);
and and303(ip_9_15,x[9],y[15]);
and and304(ip_9_16,x[9],y[16]);
and and305(ip_9_17,x[9],y[17]);
and and306(ip_9_18,x[9],y[18]);
and and307(ip_9_19,x[9],y[19]);
and and308(ip_9_20,x[9],y[20]);
and and309(ip_9_21,x[9],y[21]);
and and310(ip_9_22,x[9],y[22]);
and and311(ip_9_23,x[9],y[23]);
and and312(ip_9_24,x[9],y[24]);
and and313(ip_9_25,x[9],y[25]);
and and314(ip_9_26,x[9],y[26]);
and and315(ip_9_27,x[9],y[27]);
and and316(ip_9_28,x[9],y[28]);
and and317(ip_9_29,x[9],y[29]);
and and318(ip_9_30,x[9],y[30]);
and and319(ip_9_31,x[9],y[31]);
and and320(ip_10_0,x[10],y[0]);
and and321(ip_10_1,x[10],y[1]);
and and322(ip_10_2,x[10],y[2]);
and and323(ip_10_3,x[10],y[3]);
and and324(ip_10_4,x[10],y[4]);
and and325(ip_10_5,x[10],y[5]);
and and326(ip_10_6,x[10],y[6]);
and and327(ip_10_7,x[10],y[7]);
and and328(ip_10_8,x[10],y[8]);
and and329(ip_10_9,x[10],y[9]);
and and330(ip_10_10,x[10],y[10]);
and and331(ip_10_11,x[10],y[11]);
and and332(ip_10_12,x[10],y[12]);
and and333(ip_10_13,x[10],y[13]);
and and334(ip_10_14,x[10],y[14]);
and and335(ip_10_15,x[10],y[15]);
and and336(ip_10_16,x[10],y[16]);
and and337(ip_10_17,x[10],y[17]);
and and338(ip_10_18,x[10],y[18]);
and and339(ip_10_19,x[10],y[19]);
and and340(ip_10_20,x[10],y[20]);
and and341(ip_10_21,x[10],y[21]);
and and342(ip_10_22,x[10],y[22]);
and and343(ip_10_23,x[10],y[23]);
and and344(ip_10_24,x[10],y[24]);
and and345(ip_10_25,x[10],y[25]);
and and346(ip_10_26,x[10],y[26]);
and and347(ip_10_27,x[10],y[27]);
and and348(ip_10_28,x[10],y[28]);
and and349(ip_10_29,x[10],y[29]);
and and350(ip_10_30,x[10],y[30]);
and and351(ip_10_31,x[10],y[31]);
and and352(ip_11_0,x[11],y[0]);
and and353(ip_11_1,x[11],y[1]);
and and354(ip_11_2,x[11],y[2]);
and and355(ip_11_3,x[11],y[3]);
and and356(ip_11_4,x[11],y[4]);
and and357(ip_11_5,x[11],y[5]);
and and358(ip_11_6,x[11],y[6]);
and and359(ip_11_7,x[11],y[7]);
and and360(ip_11_8,x[11],y[8]);
and and361(ip_11_9,x[11],y[9]);
and and362(ip_11_10,x[11],y[10]);
and and363(ip_11_11,x[11],y[11]);
and and364(ip_11_12,x[11],y[12]);
and and365(ip_11_13,x[11],y[13]);
and and366(ip_11_14,x[11],y[14]);
and and367(ip_11_15,x[11],y[15]);
and and368(ip_11_16,x[11],y[16]);
and and369(ip_11_17,x[11],y[17]);
and and370(ip_11_18,x[11],y[18]);
and and371(ip_11_19,x[11],y[19]);
and and372(ip_11_20,x[11],y[20]);
and and373(ip_11_21,x[11],y[21]);
and and374(ip_11_22,x[11],y[22]);
and and375(ip_11_23,x[11],y[23]);
and and376(ip_11_24,x[11],y[24]);
and and377(ip_11_25,x[11],y[25]);
and and378(ip_11_26,x[11],y[26]);
and and379(ip_11_27,x[11],y[27]);
and and380(ip_11_28,x[11],y[28]);
and and381(ip_11_29,x[11],y[29]);
and and382(ip_11_30,x[11],y[30]);
and and383(ip_11_31,x[11],y[31]);
and and384(ip_12_0,x[12],y[0]);
and and385(ip_12_1,x[12],y[1]);
and and386(ip_12_2,x[12],y[2]);
and and387(ip_12_3,x[12],y[3]);
and and388(ip_12_4,x[12],y[4]);
and and389(ip_12_5,x[12],y[5]);
and and390(ip_12_6,x[12],y[6]);
and and391(ip_12_7,x[12],y[7]);
and and392(ip_12_8,x[12],y[8]);
and and393(ip_12_9,x[12],y[9]);
and and394(ip_12_10,x[12],y[10]);
and and395(ip_12_11,x[12],y[11]);
and and396(ip_12_12,x[12],y[12]);
and and397(ip_12_13,x[12],y[13]);
and and398(ip_12_14,x[12],y[14]);
and and399(ip_12_15,x[12],y[15]);
and and400(ip_12_16,x[12],y[16]);
and and401(ip_12_17,x[12],y[17]);
and and402(ip_12_18,x[12],y[18]);
and and403(ip_12_19,x[12],y[19]);
and and404(ip_12_20,x[12],y[20]);
and and405(ip_12_21,x[12],y[21]);
and and406(ip_12_22,x[12],y[22]);
and and407(ip_12_23,x[12],y[23]);
and and408(ip_12_24,x[12],y[24]);
and and409(ip_12_25,x[12],y[25]);
and and410(ip_12_26,x[12],y[26]);
and and411(ip_12_27,x[12],y[27]);
and and412(ip_12_28,x[12],y[28]);
and and413(ip_12_29,x[12],y[29]);
and and414(ip_12_30,x[12],y[30]);
and and415(ip_12_31,x[12],y[31]);
and and416(ip_13_0,x[13],y[0]);
and and417(ip_13_1,x[13],y[1]);
and and418(ip_13_2,x[13],y[2]);
and and419(ip_13_3,x[13],y[3]);
and and420(ip_13_4,x[13],y[4]);
and and421(ip_13_5,x[13],y[5]);
and and422(ip_13_6,x[13],y[6]);
and and423(ip_13_7,x[13],y[7]);
and and424(ip_13_8,x[13],y[8]);
and and425(ip_13_9,x[13],y[9]);
and and426(ip_13_10,x[13],y[10]);
and and427(ip_13_11,x[13],y[11]);
and and428(ip_13_12,x[13],y[12]);
and and429(ip_13_13,x[13],y[13]);
and and430(ip_13_14,x[13],y[14]);
and and431(ip_13_15,x[13],y[15]);
and and432(ip_13_16,x[13],y[16]);
and and433(ip_13_17,x[13],y[17]);
and and434(ip_13_18,x[13],y[18]);
and and435(ip_13_19,x[13],y[19]);
and and436(ip_13_20,x[13],y[20]);
and and437(ip_13_21,x[13],y[21]);
and and438(ip_13_22,x[13],y[22]);
and and439(ip_13_23,x[13],y[23]);
and and440(ip_13_24,x[13],y[24]);
and and441(ip_13_25,x[13],y[25]);
and and442(ip_13_26,x[13],y[26]);
and and443(ip_13_27,x[13],y[27]);
and and444(ip_13_28,x[13],y[28]);
and and445(ip_13_29,x[13],y[29]);
and and446(ip_13_30,x[13],y[30]);
and and447(ip_13_31,x[13],y[31]);
and and448(ip_14_0,x[14],y[0]);
and and449(ip_14_1,x[14],y[1]);
and and450(ip_14_2,x[14],y[2]);
and and451(ip_14_3,x[14],y[3]);
and and452(ip_14_4,x[14],y[4]);
and and453(ip_14_5,x[14],y[5]);
and and454(ip_14_6,x[14],y[6]);
and and455(ip_14_7,x[14],y[7]);
and and456(ip_14_8,x[14],y[8]);
and and457(ip_14_9,x[14],y[9]);
and and458(ip_14_10,x[14],y[10]);
and and459(ip_14_11,x[14],y[11]);
and and460(ip_14_12,x[14],y[12]);
and and461(ip_14_13,x[14],y[13]);
and and462(ip_14_14,x[14],y[14]);
and and463(ip_14_15,x[14],y[15]);
and and464(ip_14_16,x[14],y[16]);
and and465(ip_14_17,x[14],y[17]);
and and466(ip_14_18,x[14],y[18]);
and and467(ip_14_19,x[14],y[19]);
and and468(ip_14_20,x[14],y[20]);
and and469(ip_14_21,x[14],y[21]);
and and470(ip_14_22,x[14],y[22]);
and and471(ip_14_23,x[14],y[23]);
and and472(ip_14_24,x[14],y[24]);
and and473(ip_14_25,x[14],y[25]);
and and474(ip_14_26,x[14],y[26]);
and and475(ip_14_27,x[14],y[27]);
and and476(ip_14_28,x[14],y[28]);
and and477(ip_14_29,x[14],y[29]);
and and478(ip_14_30,x[14],y[30]);
and and479(ip_14_31,x[14],y[31]);
and and480(ip_15_0,x[15],y[0]);
and and481(ip_15_1,x[15],y[1]);
and and482(ip_15_2,x[15],y[2]);
and and483(ip_15_3,x[15],y[3]);
and and484(ip_15_4,x[15],y[4]);
and and485(ip_15_5,x[15],y[5]);
and and486(ip_15_6,x[15],y[6]);
and and487(ip_15_7,x[15],y[7]);
and and488(ip_15_8,x[15],y[8]);
and and489(ip_15_9,x[15],y[9]);
and and490(ip_15_10,x[15],y[10]);
and and491(ip_15_11,x[15],y[11]);
and and492(ip_15_12,x[15],y[12]);
and and493(ip_15_13,x[15],y[13]);
and and494(ip_15_14,x[15],y[14]);
and and495(ip_15_15,x[15],y[15]);
and and496(ip_15_16,x[15],y[16]);
and and497(ip_15_17,x[15],y[17]);
and and498(ip_15_18,x[15],y[18]);
and and499(ip_15_19,x[15],y[19]);
and and500(ip_15_20,x[15],y[20]);
and and501(ip_15_21,x[15],y[21]);
and and502(ip_15_22,x[15],y[22]);
and and503(ip_15_23,x[15],y[23]);
and and504(ip_15_24,x[15],y[24]);
and and505(ip_15_25,x[15],y[25]);
and and506(ip_15_26,x[15],y[26]);
and and507(ip_15_27,x[15],y[27]);
and and508(ip_15_28,x[15],y[28]);
and and509(ip_15_29,x[15],y[29]);
and and510(ip_15_30,x[15],y[30]);
and and511(ip_15_31,x[15],y[31]);
and and512(ip_16_0,x[16],y[0]);
and and513(ip_16_1,x[16],y[1]);
and and514(ip_16_2,x[16],y[2]);
and and515(ip_16_3,x[16],y[3]);
and and516(ip_16_4,x[16],y[4]);
and and517(ip_16_5,x[16],y[5]);
and and518(ip_16_6,x[16],y[6]);
and and519(ip_16_7,x[16],y[7]);
and and520(ip_16_8,x[16],y[8]);
and and521(ip_16_9,x[16],y[9]);
and and522(ip_16_10,x[16],y[10]);
and and523(ip_16_11,x[16],y[11]);
and and524(ip_16_12,x[16],y[12]);
and and525(ip_16_13,x[16],y[13]);
and and526(ip_16_14,x[16],y[14]);
and and527(ip_16_15,x[16],y[15]);
and and528(ip_16_16,x[16],y[16]);
and and529(ip_16_17,x[16],y[17]);
and and530(ip_16_18,x[16],y[18]);
and and531(ip_16_19,x[16],y[19]);
and and532(ip_16_20,x[16],y[20]);
and and533(ip_16_21,x[16],y[21]);
and and534(ip_16_22,x[16],y[22]);
and and535(ip_16_23,x[16],y[23]);
and and536(ip_16_24,x[16],y[24]);
and and537(ip_16_25,x[16],y[25]);
and and538(ip_16_26,x[16],y[26]);
and and539(ip_16_27,x[16],y[27]);
and and540(ip_16_28,x[16],y[28]);
and and541(ip_16_29,x[16],y[29]);
and and542(ip_16_30,x[16],y[30]);
and and543(ip_16_31,x[16],y[31]);
and and544(ip_17_0,x[17],y[0]);
and and545(ip_17_1,x[17],y[1]);
and and546(ip_17_2,x[17],y[2]);
and and547(ip_17_3,x[17],y[3]);
and and548(ip_17_4,x[17],y[4]);
and and549(ip_17_5,x[17],y[5]);
and and550(ip_17_6,x[17],y[6]);
and and551(ip_17_7,x[17],y[7]);
and and552(ip_17_8,x[17],y[8]);
and and553(ip_17_9,x[17],y[9]);
and and554(ip_17_10,x[17],y[10]);
and and555(ip_17_11,x[17],y[11]);
and and556(ip_17_12,x[17],y[12]);
and and557(ip_17_13,x[17],y[13]);
and and558(ip_17_14,x[17],y[14]);
and and559(ip_17_15,x[17],y[15]);
and and560(ip_17_16,x[17],y[16]);
and and561(ip_17_17,x[17],y[17]);
and and562(ip_17_18,x[17],y[18]);
and and563(ip_17_19,x[17],y[19]);
and and564(ip_17_20,x[17],y[20]);
and and565(ip_17_21,x[17],y[21]);
and and566(ip_17_22,x[17],y[22]);
and and567(ip_17_23,x[17],y[23]);
and and568(ip_17_24,x[17],y[24]);
and and569(ip_17_25,x[17],y[25]);
and and570(ip_17_26,x[17],y[26]);
and and571(ip_17_27,x[17],y[27]);
and and572(ip_17_28,x[17],y[28]);
and and573(ip_17_29,x[17],y[29]);
and and574(ip_17_30,x[17],y[30]);
and and575(ip_17_31,x[17],y[31]);
and and576(ip_18_0,x[18],y[0]);
and and577(ip_18_1,x[18],y[1]);
and and578(ip_18_2,x[18],y[2]);
and and579(ip_18_3,x[18],y[3]);
and and580(ip_18_4,x[18],y[4]);
and and581(ip_18_5,x[18],y[5]);
and and582(ip_18_6,x[18],y[6]);
and and583(ip_18_7,x[18],y[7]);
and and584(ip_18_8,x[18],y[8]);
and and585(ip_18_9,x[18],y[9]);
and and586(ip_18_10,x[18],y[10]);
and and587(ip_18_11,x[18],y[11]);
and and588(ip_18_12,x[18],y[12]);
and and589(ip_18_13,x[18],y[13]);
and and590(ip_18_14,x[18],y[14]);
and and591(ip_18_15,x[18],y[15]);
and and592(ip_18_16,x[18],y[16]);
and and593(ip_18_17,x[18],y[17]);
and and594(ip_18_18,x[18],y[18]);
and and595(ip_18_19,x[18],y[19]);
and and596(ip_18_20,x[18],y[20]);
and and597(ip_18_21,x[18],y[21]);
and and598(ip_18_22,x[18],y[22]);
and and599(ip_18_23,x[18],y[23]);
and and600(ip_18_24,x[18],y[24]);
and and601(ip_18_25,x[18],y[25]);
and and602(ip_18_26,x[18],y[26]);
and and603(ip_18_27,x[18],y[27]);
and and604(ip_18_28,x[18],y[28]);
and and605(ip_18_29,x[18],y[29]);
and and606(ip_18_30,x[18],y[30]);
and and607(ip_18_31,x[18],y[31]);
and and608(ip_19_0,x[19],y[0]);
and and609(ip_19_1,x[19],y[1]);
and and610(ip_19_2,x[19],y[2]);
and and611(ip_19_3,x[19],y[3]);
and and612(ip_19_4,x[19],y[4]);
and and613(ip_19_5,x[19],y[5]);
and and614(ip_19_6,x[19],y[6]);
and and615(ip_19_7,x[19],y[7]);
and and616(ip_19_8,x[19],y[8]);
and and617(ip_19_9,x[19],y[9]);
and and618(ip_19_10,x[19],y[10]);
and and619(ip_19_11,x[19],y[11]);
and and620(ip_19_12,x[19],y[12]);
and and621(ip_19_13,x[19],y[13]);
and and622(ip_19_14,x[19],y[14]);
and and623(ip_19_15,x[19],y[15]);
and and624(ip_19_16,x[19],y[16]);
and and625(ip_19_17,x[19],y[17]);
and and626(ip_19_18,x[19],y[18]);
and and627(ip_19_19,x[19],y[19]);
and and628(ip_19_20,x[19],y[20]);
and and629(ip_19_21,x[19],y[21]);
and and630(ip_19_22,x[19],y[22]);
and and631(ip_19_23,x[19],y[23]);
and and632(ip_19_24,x[19],y[24]);
and and633(ip_19_25,x[19],y[25]);
and and634(ip_19_26,x[19],y[26]);
and and635(ip_19_27,x[19],y[27]);
and and636(ip_19_28,x[19],y[28]);
and and637(ip_19_29,x[19],y[29]);
and and638(ip_19_30,x[19],y[30]);
and and639(ip_19_31,x[19],y[31]);
and and640(ip_20_0,x[20],y[0]);
and and641(ip_20_1,x[20],y[1]);
and and642(ip_20_2,x[20],y[2]);
and and643(ip_20_3,x[20],y[3]);
and and644(ip_20_4,x[20],y[4]);
and and645(ip_20_5,x[20],y[5]);
and and646(ip_20_6,x[20],y[6]);
and and647(ip_20_7,x[20],y[7]);
and and648(ip_20_8,x[20],y[8]);
and and649(ip_20_9,x[20],y[9]);
and and650(ip_20_10,x[20],y[10]);
and and651(ip_20_11,x[20],y[11]);
and and652(ip_20_12,x[20],y[12]);
and and653(ip_20_13,x[20],y[13]);
and and654(ip_20_14,x[20],y[14]);
and and655(ip_20_15,x[20],y[15]);
and and656(ip_20_16,x[20],y[16]);
and and657(ip_20_17,x[20],y[17]);
and and658(ip_20_18,x[20],y[18]);
and and659(ip_20_19,x[20],y[19]);
and and660(ip_20_20,x[20],y[20]);
and and661(ip_20_21,x[20],y[21]);
and and662(ip_20_22,x[20],y[22]);
and and663(ip_20_23,x[20],y[23]);
and and664(ip_20_24,x[20],y[24]);
and and665(ip_20_25,x[20],y[25]);
and and666(ip_20_26,x[20],y[26]);
and and667(ip_20_27,x[20],y[27]);
and and668(ip_20_28,x[20],y[28]);
and and669(ip_20_29,x[20],y[29]);
and and670(ip_20_30,x[20],y[30]);
and and671(ip_20_31,x[20],y[31]);
and and672(ip_21_0,x[21],y[0]);
and and673(ip_21_1,x[21],y[1]);
and and674(ip_21_2,x[21],y[2]);
and and675(ip_21_3,x[21],y[3]);
and and676(ip_21_4,x[21],y[4]);
and and677(ip_21_5,x[21],y[5]);
and and678(ip_21_6,x[21],y[6]);
and and679(ip_21_7,x[21],y[7]);
and and680(ip_21_8,x[21],y[8]);
and and681(ip_21_9,x[21],y[9]);
and and682(ip_21_10,x[21],y[10]);
and and683(ip_21_11,x[21],y[11]);
and and684(ip_21_12,x[21],y[12]);
and and685(ip_21_13,x[21],y[13]);
and and686(ip_21_14,x[21],y[14]);
and and687(ip_21_15,x[21],y[15]);
and and688(ip_21_16,x[21],y[16]);
and and689(ip_21_17,x[21],y[17]);
and and690(ip_21_18,x[21],y[18]);
and and691(ip_21_19,x[21],y[19]);
and and692(ip_21_20,x[21],y[20]);
and and693(ip_21_21,x[21],y[21]);
and and694(ip_21_22,x[21],y[22]);
and and695(ip_21_23,x[21],y[23]);
and and696(ip_21_24,x[21],y[24]);
and and697(ip_21_25,x[21],y[25]);
and and698(ip_21_26,x[21],y[26]);
and and699(ip_21_27,x[21],y[27]);
and and700(ip_21_28,x[21],y[28]);
and and701(ip_21_29,x[21],y[29]);
and and702(ip_21_30,x[21],y[30]);
and and703(ip_21_31,x[21],y[31]);
and and704(ip_22_0,x[22],y[0]);
and and705(ip_22_1,x[22],y[1]);
and and706(ip_22_2,x[22],y[2]);
and and707(ip_22_3,x[22],y[3]);
and and708(ip_22_4,x[22],y[4]);
and and709(ip_22_5,x[22],y[5]);
and and710(ip_22_6,x[22],y[6]);
and and711(ip_22_7,x[22],y[7]);
and and712(ip_22_8,x[22],y[8]);
and and713(ip_22_9,x[22],y[9]);
and and714(ip_22_10,x[22],y[10]);
and and715(ip_22_11,x[22],y[11]);
and and716(ip_22_12,x[22],y[12]);
and and717(ip_22_13,x[22],y[13]);
and and718(ip_22_14,x[22],y[14]);
and and719(ip_22_15,x[22],y[15]);
and and720(ip_22_16,x[22],y[16]);
and and721(ip_22_17,x[22],y[17]);
and and722(ip_22_18,x[22],y[18]);
and and723(ip_22_19,x[22],y[19]);
and and724(ip_22_20,x[22],y[20]);
and and725(ip_22_21,x[22],y[21]);
and and726(ip_22_22,x[22],y[22]);
and and727(ip_22_23,x[22],y[23]);
and and728(ip_22_24,x[22],y[24]);
and and729(ip_22_25,x[22],y[25]);
and and730(ip_22_26,x[22],y[26]);
and and731(ip_22_27,x[22],y[27]);
and and732(ip_22_28,x[22],y[28]);
and and733(ip_22_29,x[22],y[29]);
and and734(ip_22_30,x[22],y[30]);
and and735(ip_22_31,x[22],y[31]);
and and736(ip_23_0,x[23],y[0]);
and and737(ip_23_1,x[23],y[1]);
and and738(ip_23_2,x[23],y[2]);
and and739(ip_23_3,x[23],y[3]);
and and740(ip_23_4,x[23],y[4]);
and and741(ip_23_5,x[23],y[5]);
and and742(ip_23_6,x[23],y[6]);
and and743(ip_23_7,x[23],y[7]);
and and744(ip_23_8,x[23],y[8]);
and and745(ip_23_9,x[23],y[9]);
and and746(ip_23_10,x[23],y[10]);
and and747(ip_23_11,x[23],y[11]);
and and748(ip_23_12,x[23],y[12]);
and and749(ip_23_13,x[23],y[13]);
and and750(ip_23_14,x[23],y[14]);
and and751(ip_23_15,x[23],y[15]);
and and752(ip_23_16,x[23],y[16]);
and and753(ip_23_17,x[23],y[17]);
and and754(ip_23_18,x[23],y[18]);
and and755(ip_23_19,x[23],y[19]);
and and756(ip_23_20,x[23],y[20]);
and and757(ip_23_21,x[23],y[21]);
and and758(ip_23_22,x[23],y[22]);
and and759(ip_23_23,x[23],y[23]);
and and760(ip_23_24,x[23],y[24]);
and and761(ip_23_25,x[23],y[25]);
and and762(ip_23_26,x[23],y[26]);
and and763(ip_23_27,x[23],y[27]);
and and764(ip_23_28,x[23],y[28]);
and and765(ip_23_29,x[23],y[29]);
and and766(ip_23_30,x[23],y[30]);
and and767(ip_23_31,x[23],y[31]);
and and768(ip_24_0,x[24],y[0]);
and and769(ip_24_1,x[24],y[1]);
and and770(ip_24_2,x[24],y[2]);
and and771(ip_24_3,x[24],y[3]);
and and772(ip_24_4,x[24],y[4]);
and and773(ip_24_5,x[24],y[5]);
and and774(ip_24_6,x[24],y[6]);
and and775(ip_24_7,x[24],y[7]);
and and776(ip_24_8,x[24],y[8]);
and and777(ip_24_9,x[24],y[9]);
and and778(ip_24_10,x[24],y[10]);
and and779(ip_24_11,x[24],y[11]);
and and780(ip_24_12,x[24],y[12]);
and and781(ip_24_13,x[24],y[13]);
and and782(ip_24_14,x[24],y[14]);
and and783(ip_24_15,x[24],y[15]);
and and784(ip_24_16,x[24],y[16]);
and and785(ip_24_17,x[24],y[17]);
and and786(ip_24_18,x[24],y[18]);
and and787(ip_24_19,x[24],y[19]);
and and788(ip_24_20,x[24],y[20]);
and and789(ip_24_21,x[24],y[21]);
and and790(ip_24_22,x[24],y[22]);
and and791(ip_24_23,x[24],y[23]);
and and792(ip_24_24,x[24],y[24]);
and and793(ip_24_25,x[24],y[25]);
and and794(ip_24_26,x[24],y[26]);
and and795(ip_24_27,x[24],y[27]);
and and796(ip_24_28,x[24],y[28]);
and and797(ip_24_29,x[24],y[29]);
and and798(ip_24_30,x[24],y[30]);
and and799(ip_24_31,x[24],y[31]);
and and800(ip_25_0,x[25],y[0]);
and and801(ip_25_1,x[25],y[1]);
and and802(ip_25_2,x[25],y[2]);
and and803(ip_25_3,x[25],y[3]);
and and804(ip_25_4,x[25],y[4]);
and and805(ip_25_5,x[25],y[5]);
and and806(ip_25_6,x[25],y[6]);
and and807(ip_25_7,x[25],y[7]);
and and808(ip_25_8,x[25],y[8]);
and and809(ip_25_9,x[25],y[9]);
and and810(ip_25_10,x[25],y[10]);
and and811(ip_25_11,x[25],y[11]);
and and812(ip_25_12,x[25],y[12]);
and and813(ip_25_13,x[25],y[13]);
and and814(ip_25_14,x[25],y[14]);
and and815(ip_25_15,x[25],y[15]);
and and816(ip_25_16,x[25],y[16]);
and and817(ip_25_17,x[25],y[17]);
and and818(ip_25_18,x[25],y[18]);
and and819(ip_25_19,x[25],y[19]);
and and820(ip_25_20,x[25],y[20]);
and and821(ip_25_21,x[25],y[21]);
and and822(ip_25_22,x[25],y[22]);
and and823(ip_25_23,x[25],y[23]);
and and824(ip_25_24,x[25],y[24]);
and and825(ip_25_25,x[25],y[25]);
and and826(ip_25_26,x[25],y[26]);
and and827(ip_25_27,x[25],y[27]);
and and828(ip_25_28,x[25],y[28]);
and and829(ip_25_29,x[25],y[29]);
and and830(ip_25_30,x[25],y[30]);
and and831(ip_25_31,x[25],y[31]);
and and832(ip_26_0,x[26],y[0]);
and and833(ip_26_1,x[26],y[1]);
and and834(ip_26_2,x[26],y[2]);
and and835(ip_26_3,x[26],y[3]);
and and836(ip_26_4,x[26],y[4]);
and and837(ip_26_5,x[26],y[5]);
and and838(ip_26_6,x[26],y[6]);
and and839(ip_26_7,x[26],y[7]);
and and840(ip_26_8,x[26],y[8]);
and and841(ip_26_9,x[26],y[9]);
and and842(ip_26_10,x[26],y[10]);
and and843(ip_26_11,x[26],y[11]);
and and844(ip_26_12,x[26],y[12]);
and and845(ip_26_13,x[26],y[13]);
and and846(ip_26_14,x[26],y[14]);
and and847(ip_26_15,x[26],y[15]);
and and848(ip_26_16,x[26],y[16]);
and and849(ip_26_17,x[26],y[17]);
and and850(ip_26_18,x[26],y[18]);
and and851(ip_26_19,x[26],y[19]);
and and852(ip_26_20,x[26],y[20]);
and and853(ip_26_21,x[26],y[21]);
and and854(ip_26_22,x[26],y[22]);
and and855(ip_26_23,x[26],y[23]);
and and856(ip_26_24,x[26],y[24]);
and and857(ip_26_25,x[26],y[25]);
and and858(ip_26_26,x[26],y[26]);
and and859(ip_26_27,x[26],y[27]);
and and860(ip_26_28,x[26],y[28]);
and and861(ip_26_29,x[26],y[29]);
and and862(ip_26_30,x[26],y[30]);
and and863(ip_26_31,x[26],y[31]);
and and864(ip_27_0,x[27],y[0]);
and and865(ip_27_1,x[27],y[1]);
and and866(ip_27_2,x[27],y[2]);
and and867(ip_27_3,x[27],y[3]);
and and868(ip_27_4,x[27],y[4]);
and and869(ip_27_5,x[27],y[5]);
and and870(ip_27_6,x[27],y[6]);
and and871(ip_27_7,x[27],y[7]);
and and872(ip_27_8,x[27],y[8]);
and and873(ip_27_9,x[27],y[9]);
and and874(ip_27_10,x[27],y[10]);
and and875(ip_27_11,x[27],y[11]);
and and876(ip_27_12,x[27],y[12]);
and and877(ip_27_13,x[27],y[13]);
and and878(ip_27_14,x[27],y[14]);
and and879(ip_27_15,x[27],y[15]);
and and880(ip_27_16,x[27],y[16]);
and and881(ip_27_17,x[27],y[17]);
and and882(ip_27_18,x[27],y[18]);
and and883(ip_27_19,x[27],y[19]);
and and884(ip_27_20,x[27],y[20]);
and and885(ip_27_21,x[27],y[21]);
and and886(ip_27_22,x[27],y[22]);
and and887(ip_27_23,x[27],y[23]);
and and888(ip_27_24,x[27],y[24]);
and and889(ip_27_25,x[27],y[25]);
and and890(ip_27_26,x[27],y[26]);
and and891(ip_27_27,x[27],y[27]);
and and892(ip_27_28,x[27],y[28]);
and and893(ip_27_29,x[27],y[29]);
and and894(ip_27_30,x[27],y[30]);
and and895(ip_27_31,x[27],y[31]);
and and896(ip_28_0,x[28],y[0]);
and and897(ip_28_1,x[28],y[1]);
and and898(ip_28_2,x[28],y[2]);
and and899(ip_28_3,x[28],y[3]);
and and900(ip_28_4,x[28],y[4]);
and and901(ip_28_5,x[28],y[5]);
and and902(ip_28_6,x[28],y[6]);
and and903(ip_28_7,x[28],y[7]);
and and904(ip_28_8,x[28],y[8]);
and and905(ip_28_9,x[28],y[9]);
and and906(ip_28_10,x[28],y[10]);
and and907(ip_28_11,x[28],y[11]);
and and908(ip_28_12,x[28],y[12]);
and and909(ip_28_13,x[28],y[13]);
and and910(ip_28_14,x[28],y[14]);
and and911(ip_28_15,x[28],y[15]);
and and912(ip_28_16,x[28],y[16]);
and and913(ip_28_17,x[28],y[17]);
and and914(ip_28_18,x[28],y[18]);
and and915(ip_28_19,x[28],y[19]);
and and916(ip_28_20,x[28],y[20]);
and and917(ip_28_21,x[28],y[21]);
and and918(ip_28_22,x[28],y[22]);
and and919(ip_28_23,x[28],y[23]);
and and920(ip_28_24,x[28],y[24]);
and and921(ip_28_25,x[28],y[25]);
and and922(ip_28_26,x[28],y[26]);
and and923(ip_28_27,x[28],y[27]);
and and924(ip_28_28,x[28],y[28]);
and and925(ip_28_29,x[28],y[29]);
and and926(ip_28_30,x[28],y[30]);
and and927(ip_28_31,x[28],y[31]);
and and928(ip_29_0,x[29],y[0]);
and and929(ip_29_1,x[29],y[1]);
and and930(ip_29_2,x[29],y[2]);
and and931(ip_29_3,x[29],y[3]);
and and932(ip_29_4,x[29],y[4]);
and and933(ip_29_5,x[29],y[5]);
and and934(ip_29_6,x[29],y[6]);
and and935(ip_29_7,x[29],y[7]);
and and936(ip_29_8,x[29],y[8]);
and and937(ip_29_9,x[29],y[9]);
and and938(ip_29_10,x[29],y[10]);
and and939(ip_29_11,x[29],y[11]);
and and940(ip_29_12,x[29],y[12]);
and and941(ip_29_13,x[29],y[13]);
and and942(ip_29_14,x[29],y[14]);
and and943(ip_29_15,x[29],y[15]);
and and944(ip_29_16,x[29],y[16]);
and and945(ip_29_17,x[29],y[17]);
and and946(ip_29_18,x[29],y[18]);
and and947(ip_29_19,x[29],y[19]);
and and948(ip_29_20,x[29],y[20]);
and and949(ip_29_21,x[29],y[21]);
and and950(ip_29_22,x[29],y[22]);
and and951(ip_29_23,x[29],y[23]);
and and952(ip_29_24,x[29],y[24]);
and and953(ip_29_25,x[29],y[25]);
and and954(ip_29_26,x[29],y[26]);
and and955(ip_29_27,x[29],y[27]);
and and956(ip_29_28,x[29],y[28]);
and and957(ip_29_29,x[29],y[29]);
and and958(ip_29_30,x[29],y[30]);
and and959(ip_29_31,x[29],y[31]);
and and960(ip_30_0,x[30],y[0]);
and and961(ip_30_1,x[30],y[1]);
and and962(ip_30_2,x[30],y[2]);
and and963(ip_30_3,x[30],y[3]);
and and964(ip_30_4,x[30],y[4]);
and and965(ip_30_5,x[30],y[5]);
and and966(ip_30_6,x[30],y[6]);
and and967(ip_30_7,x[30],y[7]);
and and968(ip_30_8,x[30],y[8]);
and and969(ip_30_9,x[30],y[9]);
and and970(ip_30_10,x[30],y[10]);
and and971(ip_30_11,x[30],y[11]);
and and972(ip_30_12,x[30],y[12]);
and and973(ip_30_13,x[30],y[13]);
and and974(ip_30_14,x[30],y[14]);
and and975(ip_30_15,x[30],y[15]);
and and976(ip_30_16,x[30],y[16]);
and and977(ip_30_17,x[30],y[17]);
and and978(ip_30_18,x[30],y[18]);
and and979(ip_30_19,x[30],y[19]);
and and980(ip_30_20,x[30],y[20]);
and and981(ip_30_21,x[30],y[21]);
and and982(ip_30_22,x[30],y[22]);
and and983(ip_30_23,x[30],y[23]);
and and984(ip_30_24,x[30],y[24]);
and and985(ip_30_25,x[30],y[25]);
and and986(ip_30_26,x[30],y[26]);
and and987(ip_30_27,x[30],y[27]);
and and988(ip_30_28,x[30],y[28]);
and and989(ip_30_29,x[30],y[29]);
and and990(ip_30_30,x[30],y[30]);
and and991(ip_30_31,x[30],y[31]);
and and992(ip_31_0,x[31],y[0]);
and and993(ip_31_1,x[31],y[1]);
and and994(ip_31_2,x[31],y[2]);
and and995(ip_31_3,x[31],y[3]);
and and996(ip_31_4,x[31],y[4]);
and and997(ip_31_5,x[31],y[5]);
and and998(ip_31_6,x[31],y[6]);
and and999(ip_31_7,x[31],y[7]);
and and1000(ip_31_8,x[31],y[8]);
and and1001(ip_31_9,x[31],y[9]);
and and1002(ip_31_10,x[31],y[10]);
and and1003(ip_31_11,x[31],y[11]);
and and1004(ip_31_12,x[31],y[12]);
and and1005(ip_31_13,x[31],y[13]);
and and1006(ip_31_14,x[31],y[14]);
and and1007(ip_31_15,x[31],y[15]);
and and1008(ip_31_16,x[31],y[16]);
and and1009(ip_31_17,x[31],y[17]);
and and1010(ip_31_18,x[31],y[18]);
and and1011(ip_31_19,x[31],y[19]);
and and1012(ip_31_20,x[31],y[20]);
and and1013(ip_31_21,x[31],y[21]);
and and1014(ip_31_22,x[31],y[22]);
and and1015(ip_31_23,x[31],y[23]);
and and1016(ip_31_24,x[31],y[24]);
and and1017(ip_31_25,x[31],y[25]);
and and1018(ip_31_26,x[31],y[26]);
and and1019(ip_31_27,x[31],y[27]);
and and1020(ip_31_28,x[31],y[28]);
and and1021(ip_31_29,x[31],y[29]);
and and1022(ip_31_30,x[31],y[30]);
and and1023(ip_31_31,x[31],y[31]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
FA fa2(ip_3_0,p3,p0,p4,p5);
FA fa3(ip_0_4,ip_1_3,ip_2_2,p6,p7);
FA fa4(ip_3_1,ip_4_0,p7,p8,p9);
FA fa5(p2,p9,p4,p10,p11);
FA fa6(ip_0_5,ip_1_4,ip_2_3,p12,p13);
FA fa7(ip_3_2,ip_4_1,ip_5_0,p14,p15);
FA fa8(p13,p15,p6,p16,p17);
FA fa9(p17,p8,p10,p18,p19);
FA fa10(ip_0_6,ip_1_5,ip_2_4,p20,p21);
FA fa11(ip_3_3,ip_4_2,ip_5_1,p22,p23);
FA fa12(ip_6_0,p21,p23,p24,p25);
FA fa13(p12,p14,p25,p26,p27);
FA fa14(p16,p27,p18,p28,p29);
FA fa15(ip_0_7,ip_1_6,ip_2_5,p30,p31);
FA fa16(ip_3_4,ip_4_3,ip_5_2,p32,p33);
FA fa17(ip_6_1,ip_7_0,p31,p34,p35);
FA fa18(p33,p20,p22,p36,p37);
FA fa19(p35,p24,p37,p38,p39);
HA ha0(p26,p39,p40,p41);
FA fa20(ip_0_8,ip_1_7,ip_2_6,p42,p43);
FA fa21(ip_3_5,ip_4_4,ip_5_3,p44,p45);
FA fa22(ip_6_2,ip_7_1,ip_8_0,p46,p47);
FA fa23(p43,p45,p47,p48,p49);
FA fa24(p30,p32,p34,p50,p51);
FA fa25(p49,p51,p36,p52,p53);
FA fa26(p53,p38,p40,p54,p55);
FA fa27(ip_0_9,ip_1_8,ip_2_7,p56,p57);
FA fa28(ip_3_6,ip_4_5,ip_5_4,p58,p59);
FA fa29(ip_6_3,ip_7_2,ip_8_1,p60,p61);
FA fa30(ip_9_0,p57,p59,p62,p63);
FA fa31(p61,p42,p44,p64,p65);
FA fa32(p46,p63,p48,p66,p67);
FA fa33(p65,p50,p67,p68,p69);
FA fa34(p52,p69,p54,p70,p71);
FA fa35(ip_0_10,ip_1_9,ip_2_8,p72,p73);
FA fa36(ip_3_7,ip_4_6,ip_5_5,p74,p75);
FA fa37(ip_6_4,ip_7_3,ip_8_2,p76,p77);
FA fa38(ip_9_1,ip_10_0,p73,p78,p79);
FA fa39(p75,p77,p56,p80,p81);
HA ha1(p58,p60,p82,p83);
FA fa40(p79,p81,p83,p84,p85);
FA fa41(p62,p64,p85,p86,p87);
FA fa42(p66,p87,p68,p88,p89);
FA fa43(ip_0_11,ip_1_10,ip_2_9,p90,p91);
FA fa44(ip_3_8,ip_4_7,ip_5_6,p92,p93);
FA fa45(ip_6_5,ip_7_4,ip_8_3,p94,p95);
FA fa46(ip_9_2,ip_10_1,ip_11_0,p96,p97);
FA fa47(p91,p93,p95,p98,p99);
FA fa48(p97,p72,p74,p100,p101);
FA fa49(p76,p78,p82,p102,p103);
FA fa50(p99,p101,p80,p104,p105);
FA fa51(p103,p105,p84,p106,p107);
HA ha2(p107,p86,p108,p109);
FA fa52(ip_0_12,ip_1_11,ip_2_10,p110,p111);
FA fa53(ip_3_9,ip_4_8,ip_5_7,p112,p113);
FA fa54(ip_6_6,ip_7_5,ip_8_4,p114,p115);
FA fa55(ip_9_3,ip_10_2,ip_11_1,p116,p117);
FA fa56(ip_12_0,p111,p113,p118,p119);
FA fa57(p115,p117,p90,p120,p121);
FA fa58(p92,p94,p96,p122,p123);
FA fa59(p119,p121,p123,p124,p125);
FA fa60(p98,p100,p125,p126,p127);
HA ha3(p102,p104,p128,p129);
FA fa61(p127,p129,p106,p130,p131);
FA fa62(ip_0_13,ip_1_12,ip_2_11,p132,p133);
FA fa63(ip_3_10,ip_4_9,ip_5_8,p134,p135);
FA fa64(ip_6_7,ip_7_6,ip_8_5,p136,p137);
FA fa65(ip_9_4,ip_10_3,ip_11_2,p138,p139);
FA fa66(ip_12_1,ip_13_0,p133,p140,p141);
HA ha4(p135,p137,p142,p143);
FA fa67(p139,p110,p112,p144,p145);
FA fa68(p114,p116,p141,p146,p147);
FA fa69(p143,p118,p120,p148,p149);
FA fa70(p145,p147,p122,p150,p151);
FA fa71(p124,p149,p151,p152,p153);
FA fa72(p126,p128,p153,p154,p155);
FA fa73(ip_0_14,ip_1_13,ip_2_12,p156,p157);
FA fa74(ip_3_11,ip_4_10,ip_5_9,p158,p159);
FA fa75(ip_6_8,ip_7_7,ip_8_6,p160,p161);
FA fa76(ip_9_5,ip_10_4,ip_11_3,p162,p163);
FA fa77(ip_12_2,ip_13_1,ip_14_0,p164,p165);
FA fa78(p157,p159,p161,p166,p167);
FA fa79(p163,p165,p132,p168,p169);
FA fa80(p134,p136,p138,p170,p171);
FA fa81(p142,p140,p167,p172,p173);
FA fa82(p169,p171,p144,p174,p175);
HA ha5(p146,p173,p176,p177);
FA fa83(p175,p177,p148,p178,p179);
FA fa84(p150,p179,p152,p180,p181);
FA fa85(ip_0_15,ip_1_14,ip_2_13,p182,p183);
HA ha6(ip_3_12,ip_4_11,p184,p185);
FA fa86(ip_5_10,ip_6_9,ip_7_8,p186,p187);
FA fa87(ip_8_7,ip_9_6,ip_10_5,p188,p189);
HA ha7(ip_11_4,ip_12_3,p190,p191);
FA fa88(ip_13_2,ip_14_1,ip_15_0,p192,p193);
FA fa89(p185,p191,p183,p194,p195);
FA fa90(p187,p189,p193,p196,p197);
FA fa91(p156,p158,p160,p198,p199);
FA fa92(p162,p164,p195,p200,p201);
FA fa93(p197,p166,p168,p202,p203);
FA fa94(p199,p201,p170,p204,p205);
HA ha8(p172,p176,p206,p207);
FA fa95(p203,p205,p174,p208,p209);
FA fa96(p207,p209,p178,p210,p211);
HA ha9(ip_0_16,ip_1_15,p212,p213);
FA fa97(ip_2_14,ip_3_13,ip_4_12,p214,p215);
FA fa98(ip_5_11,ip_6_10,ip_7_9,p216,p217);
FA fa99(ip_8_8,ip_9_7,ip_10_6,p218,p219);
FA fa100(ip_11_5,ip_12_4,ip_13_3,p220,p221);
FA fa101(ip_14_2,ip_15_1,ip_16_0,p222,p223);
FA fa102(p184,p190,p213,p224,p225);
FA fa103(p215,p217,p219,p226,p227);
FA fa104(p221,p223,p182,p228,p229);
FA fa105(p186,p188,p192,p230,p231);
FA fa106(p225,p194,p227,p232,p233);
FA fa107(p229,p196,p231,p234,p235);
FA fa108(p198,p200,p233,p236,p237);
FA fa109(p235,p202,p204,p238,p239);
FA fa110(p206,p237,p208,p240,p241);
FA fa111(p239,p241,p210,p242,p243);
HA ha10(ip_0_17,ip_1_16,p244,p245);
FA fa112(ip_2_15,ip_3_14,ip_4_13,p246,p247);
FA fa113(ip_5_12,ip_6_11,ip_7_10,p248,p249);
FA fa114(ip_8_9,ip_9_8,ip_10_7,p250,p251);
FA fa115(ip_11_6,ip_12_5,ip_13_4,p252,p253);
FA fa116(ip_14_3,ip_15_2,ip_16_1,p254,p255);
FA fa117(ip_17_0,p212,p245,p256,p257);
FA fa118(p247,p249,p251,p258,p259);
FA fa119(p253,p255,p214,p260,p261);
FA fa120(p216,p218,p220,p262,p263);
FA fa121(p222,p257,p224,p264,p265);
FA fa122(p259,p261,p226,p266,p267);
FA fa123(p228,p263,p265,p268,p269);
FA fa124(p230,p267,p232,p270,p271);
FA fa125(p269,p234,p271,p272,p273);
FA fa126(p236,p273,p238,p274,p275);
FA fa127(p240,p275,p242,p276,p277);
FA fa128(ip_0_18,ip_1_17,ip_2_16,p278,p279);
FA fa129(ip_3_15,ip_4_14,ip_5_13,p280,p281);
FA fa130(ip_6_12,ip_7_11,ip_8_10,p282,p283);
FA fa131(ip_9_9,ip_10_8,ip_11_7,p284,p285);
FA fa132(ip_12_6,ip_13_5,ip_14_4,p286,p287);
FA fa133(ip_15_3,ip_16_2,ip_17_1,p288,p289);
FA fa134(ip_18_0,p244,p279,p290,p291);
FA fa135(p281,p283,p285,p292,p293);
FA fa136(p287,p289,p246,p294,p295);
FA fa137(p248,p250,p252,p296,p297);
FA fa138(p254,p291,p256,p298,p299);
FA fa139(p293,p295,p258,p300,p301);
FA fa140(p260,p297,p299,p302,p303);
FA fa141(p262,p264,p301,p304,p305);
FA fa142(p266,p303,p268,p306,p307);
FA fa143(p305,p270,p307,p308,p309);
FA fa144(p272,p309,p274,p310,p311);
FA fa145(ip_0_19,ip_1_18,ip_2_17,p312,p313);
FA fa146(ip_3_16,ip_4_15,ip_5_14,p314,p315);
FA fa147(ip_6_13,ip_7_12,ip_8_11,p316,p317);
FA fa148(ip_9_10,ip_10_9,ip_11_8,p318,p319);
FA fa149(ip_12_7,ip_13_6,ip_14_5,p320,p321);
FA fa150(ip_15_4,ip_16_3,ip_17_2,p322,p323);
FA fa151(ip_18_1,ip_19_0,p313,p324,p325);
FA fa152(p315,p317,p319,p326,p327);
FA fa153(p321,p323,p278,p328,p329);
FA fa154(p280,p282,p284,p330,p331);
FA fa155(p286,p288,p325,p332,p333);
FA fa156(p290,p327,p329,p334,p335);
HA ha11(p292,p294,p336,p337);
FA fa157(p331,p333,p296,p338,p339);
FA fa158(p298,p335,p337,p340,p341);
FA fa159(p300,p339,p302,p342,p343);
FA fa160(p341,p304,p343,p344,p345);
HA ha12(p306,p345,p346,p347);
FA fa161(p308,p347,p310,p348,p349);
FA fa162(ip_0_20,ip_1_19,ip_2_18,p350,p351);
FA fa163(ip_3_17,ip_4_16,ip_5_15,p352,p353);
FA fa164(ip_6_14,ip_7_13,ip_8_12,p354,p355);
FA fa165(ip_9_11,ip_10_10,ip_11_9,p356,p357);
FA fa166(ip_12_8,ip_13_7,ip_14_6,p358,p359);
HA ha13(ip_15_5,ip_16_4,p360,p361);
FA fa167(ip_17_3,ip_18_2,ip_19_1,p362,p363);
FA fa168(ip_20_0,p361,p351,p364,p365);
FA fa169(p353,p355,p357,p366,p367);
FA fa170(p359,p363,p312,p368,p369);
FA fa171(p314,p316,p318,p370,p371);
FA fa172(p320,p322,p365,p372,p373);
FA fa173(p324,p367,p369,p374,p375);
FA fa174(p326,p328,p371,p376,p377);
FA fa175(p373,p330,p332,p378,p379);
FA fa176(p336,p375,p334,p380,p381);
FA fa177(p377,p338,p379,p382,p383);
FA fa178(p381,p340,p342,p384,p385);
FA fa179(p383,p385,p344,p386,p387);
FA fa180(p346,p387,p348,p388,p389);
FA fa181(ip_0_21,ip_1_20,ip_2_19,p390,p391);
FA fa182(ip_3_18,ip_4_17,ip_5_16,p392,p393);
FA fa183(ip_6_15,ip_7_14,ip_8_13,p394,p395);
FA fa184(ip_9_12,ip_10_11,ip_11_10,p396,p397);
FA fa185(ip_12_9,ip_13_8,ip_14_7,p398,p399);
FA fa186(ip_15_6,ip_16_5,ip_17_4,p400,p401);
FA fa187(ip_18_3,ip_19_2,ip_20_1,p402,p403);
FA fa188(ip_21_0,p360,p391,p404,p405);
FA fa189(p393,p395,p397,p406,p407);
FA fa190(p399,p401,p403,p408,p409);
FA fa191(p350,p352,p354,p410,p411);
FA fa192(p356,p358,p362,p412,p413);
FA fa193(p405,p364,p407,p414,p415);
FA fa194(p409,p366,p368,p416,p417);
FA fa195(p411,p413,p370,p418,p419);
FA fa196(p372,p415,p374,p420,p421);
FA fa197(p417,p419,p376,p422,p423);
FA fa198(p421,p378,p380,p424,p425);
FA fa199(p423,p382,p425,p426,p427);
FA fa200(p384,p427,p386,p428,p429);
FA fa201(ip_0_22,ip_1_21,ip_2_20,p430,p431);
FA fa202(ip_3_19,ip_4_18,ip_5_17,p432,p433);
FA fa203(ip_6_16,ip_7_15,ip_8_14,p434,p435);
FA fa204(ip_9_13,ip_10_12,ip_11_11,p436,p437);
FA fa205(ip_12_10,ip_13_9,ip_14_8,p438,p439);
FA fa206(ip_15_7,ip_16_6,ip_17_5,p440,p441);
FA fa207(ip_18_4,ip_19_3,ip_20_2,p442,p443);
FA fa208(ip_21_1,ip_22_0,p431,p444,p445);
FA fa209(p433,p435,p437,p446,p447);
FA fa210(p439,p441,p443,p448,p449);
FA fa211(p390,p392,p394,p450,p451);
FA fa212(p396,p398,p400,p452,p453);
FA fa213(p402,p445,p404,p454,p455);
FA fa214(p447,p449,p406,p456,p457);
FA fa215(p408,p451,p453,p458,p459);
FA fa216(p455,p410,p412,p460,p461);
FA fa217(p457,p414,p459,p462,p463);
FA fa218(p416,p418,p461,p464,p465);
FA fa219(p420,p463,p422,p466,p467);
FA fa220(p465,p467,p424,p468,p469);
FA fa221(p469,p426,p428,p470,p471);
FA fa222(ip_0_23,ip_1_22,ip_2_21,p472,p473);
FA fa223(ip_3_20,ip_4_19,ip_5_18,p474,p475);
FA fa224(ip_6_17,ip_7_16,ip_8_15,p476,p477);
FA fa225(ip_9_14,ip_10_13,ip_11_12,p478,p479);
FA fa226(ip_12_11,ip_13_10,ip_14_9,p480,p481);
FA fa227(ip_15_8,ip_16_7,ip_17_6,p482,p483);
FA fa228(ip_18_5,ip_19_4,ip_20_3,p484,p485);
FA fa229(ip_21_2,ip_22_1,ip_23_0,p486,p487);
FA fa230(p473,p475,p477,p488,p489);
FA fa231(p479,p481,p483,p490,p491);
FA fa232(p485,p487,p430,p492,p493);
FA fa233(p432,p434,p436,p494,p495);
FA fa234(p438,p440,p442,p496,p497);
FA fa235(p444,p489,p491,p498,p499);
FA fa236(p493,p446,p448,p500,p501);
FA fa237(p495,p497,p450,p502,p503);
FA fa238(p452,p454,p499,p504,p505);
FA fa239(p456,p501,p503,p506,p507);
FA fa240(p458,p505,p460,p508,p509);
FA fa241(p507,p462,p509,p510,p511);
FA fa242(p464,p466,p511,p512,p513);
FA fa243(p468,p513,p470,p514,p515);
FA fa244(ip_0_24,ip_1_23,ip_2_22,p516,p517);
FA fa245(ip_3_21,ip_4_20,ip_5_19,p518,p519);
FA fa246(ip_6_18,ip_7_17,ip_8_16,p520,p521);
FA fa247(ip_9_15,ip_10_14,ip_11_13,p522,p523);
FA fa248(ip_12_12,ip_13_11,ip_14_10,p524,p525);
FA fa249(ip_15_9,ip_16_8,ip_17_7,p526,p527);
FA fa250(ip_18_6,ip_19_5,ip_20_4,p528,p529);
FA fa251(ip_21_3,ip_22_2,ip_23_1,p530,p531);
FA fa252(ip_24_0,p517,p519,p532,p533);
FA fa253(p521,p523,p525,p534,p535);
HA ha14(p527,p529,p536,p537);
FA fa254(p531,p472,p474,p538,p539);
FA fa255(p476,p478,p480,p540,p541);
FA fa256(p482,p484,p486,p542,p543);
FA fa257(p537,p533,p535,p544,p545);
FA fa258(p488,p490,p492,p546,p547);
FA fa259(p539,p541,p543,p548,p549);
FA fa260(p494,p496,p545,p550,p551);
FA fa261(p498,p547,p549,p552,p553);
FA fa262(p500,p502,p551,p554,p555);
HA ha15(p504,p553,p556,p557);
FA fa263(p506,p555,p557,p558,p559);
FA fa264(p508,p559,p510,p560,p561);
HA ha16(p561,p512,p562,p563);
FA fa265(ip_0_25,ip_1_24,ip_2_23,p564,p565);
HA ha17(ip_3_22,ip_4_21,p566,p567);
FA fa266(ip_5_20,ip_6_19,ip_7_18,p568,p569);
FA fa267(ip_8_17,ip_9_16,ip_10_15,p570,p571);
FA fa268(ip_11_14,ip_12_13,ip_13_12,p572,p573);
FA fa269(ip_14_11,ip_15_10,ip_16_9,p574,p575);
FA fa270(ip_17_8,ip_18_7,ip_19_6,p576,p577);
FA fa271(ip_20_5,ip_21_4,ip_22_3,p578,p579);
FA fa272(ip_23_2,ip_24_1,ip_25_0,p580,p581);
FA fa273(p567,p565,p569,p582,p583);
FA fa274(p571,p573,p575,p584,p585);
FA fa275(p577,p579,p581,p586,p587);
FA fa276(p516,p518,p520,p588,p589);
FA fa277(p522,p524,p526,p590,p591);
FA fa278(p528,p530,p536,p592,p593);
FA fa279(p583,p585,p587,p594,p595);
FA fa280(p532,p534,p589,p596,p597);
FA fa281(p591,p593,p538,p598,p599);
FA fa282(p540,p542,p595,p600,p601);
FA fa283(p544,p597,p599,p602,p603);
FA fa284(p546,p548,p601,p604,p605);
FA fa285(p550,p603,p552,p606,p607);
FA fa286(p556,p605,p554,p608,p609);
FA fa287(p607,p609,p558,p610,p611);
FA fa288(p611,p560,p562,p612,p613);
FA fa289(ip_0_26,ip_1_25,ip_2_24,p614,p615);
HA ha18(ip_3_23,ip_4_22,p616,p617);
FA fa290(ip_5_21,ip_6_20,ip_7_19,p618,p619);
FA fa291(ip_8_18,ip_9_17,ip_10_16,p620,p621);
HA ha19(ip_11_15,ip_12_14,p622,p623);
FA fa292(ip_13_13,ip_14_12,ip_15_11,p624,p625);
FA fa293(ip_16_10,ip_17_9,ip_18_8,p626,p627);
FA fa294(ip_19_7,ip_20_6,ip_21_5,p628,p629);
FA fa295(ip_22_4,ip_23_3,ip_24_2,p630,p631);
FA fa296(ip_25_1,ip_26_0,p566,p632,p633);
FA fa297(p617,p623,p615,p634,p635);
FA fa298(p619,p621,p625,p636,p637);
FA fa299(p627,p629,p631,p638,p639);
FA fa300(p633,p564,p568,p640,p641);
FA fa301(p570,p572,p574,p642,p643);
FA fa302(p576,p578,p580,p644,p645);
FA fa303(p635,p637,p639,p646,p647);
FA fa304(p582,p584,p586,p648,p649);
FA fa305(p641,p643,p645,p650,p651);
FA fa306(p588,p590,p592,p652,p653);
FA fa307(p647,p594,p649,p654,p655);
FA fa308(p651,p596,p598,p656,p657);
FA fa309(p653,p600,p655,p658,p659);
FA fa310(p602,p657,p604,p660,p661);
FA fa311(p659,p606,p661,p662,p663);
FA fa312(p608,p663,p610,p664,p665);
FA fa313(ip_0_27,ip_1_26,ip_2_25,p666,p667);
FA fa314(ip_3_24,ip_4_23,ip_5_22,p668,p669);
FA fa315(ip_6_21,ip_7_20,ip_8_19,p670,p671);
FA fa316(ip_9_18,ip_10_17,ip_11_16,p672,p673);
FA fa317(ip_12_15,ip_13_14,ip_14_13,p674,p675);
FA fa318(ip_15_12,ip_16_11,ip_17_10,p676,p677);
FA fa319(ip_18_9,ip_19_8,ip_20_7,p678,p679);
FA fa320(ip_21_6,ip_22_5,ip_23_4,p680,p681);
FA fa321(ip_24_3,ip_25_2,ip_26_1,p682,p683);
FA fa322(ip_27_0,p616,p622,p684,p685);
FA fa323(p667,p669,p671,p686,p687);
FA fa324(p673,p675,p677,p688,p689);
FA fa325(p679,p681,p683,p690,p691);
FA fa326(p614,p618,p620,p692,p693);
FA fa327(p624,p626,p628,p694,p695);
FA fa328(p630,p632,p685,p696,p697);
FA fa329(p634,p687,p689,p698,p699);
HA ha20(p691,p636,p700,p701);
FA fa330(p638,p693,p695,p702,p703);
FA fa331(p697,p640,p642,p704,p705);
FA fa332(p644,p699,p701,p706,p707);
FA fa333(p646,p703,p648,p708,p709);
HA ha21(p650,p705,p710,p711);
FA fa334(p707,p652,p709,p712,p713);
FA fa335(p711,p654,p656,p714,p715);
FA fa336(p713,p658,p715,p716,p717);
FA fa337(p660,p717,p662,p718,p719);
FA fa338(ip_0_28,ip_1_27,ip_2_26,p720,p721);
FA fa339(ip_3_25,ip_4_24,ip_5_23,p722,p723);
FA fa340(ip_6_22,ip_7_21,ip_8_20,p724,p725);
FA fa341(ip_9_19,ip_10_18,ip_11_17,p726,p727);
FA fa342(ip_12_16,ip_13_15,ip_14_14,p728,p729);
FA fa343(ip_15_13,ip_16_12,ip_17_11,p730,p731);
FA fa344(ip_18_10,ip_19_9,ip_20_8,p732,p733);
FA fa345(ip_21_7,ip_22_6,ip_23_5,p734,p735);
FA fa346(ip_24_4,ip_25_3,ip_26_2,p736,p737);
FA fa347(ip_27_1,ip_28_0,p721,p738,p739);
HA ha22(p723,p725,p740,p741);
FA fa348(p727,p729,p731,p742,p743);
FA fa349(p733,p735,p737,p744,p745);
FA fa350(p666,p668,p670,p746,p747);
FA fa351(p672,p674,p676,p748,p749);
FA fa352(p678,p680,p682,p750,p751);
FA fa353(p739,p741,p684,p752,p753);
FA fa354(p743,p745,p686,p754,p755);
FA fa355(p688,p690,p747,p756,p757);
FA fa356(p749,p751,p753,p758,p759);
FA fa357(p692,p694,p696,p760,p761);
FA fa358(p700,p755,p698,p762,p763);
FA fa359(p757,p759,p702,p764,p765);
FA fa360(p761,p763,p704,p766,p767);
FA fa361(p706,p710,p765,p768,p769);
FA fa362(p708,p767,p769,p770,p771);
FA fa363(p712,p771,p714,p772,p773);
FA fa364(p773,p716,p718,p774,p775);
FA fa365(ip_0_29,ip_1_28,ip_2_27,p776,p777);
FA fa366(ip_3_26,ip_4_25,ip_5_24,p778,p779);
FA fa367(ip_6_23,ip_7_22,ip_8_21,p780,p781);
FA fa368(ip_9_20,ip_10_19,ip_11_18,p782,p783);
FA fa369(ip_12_17,ip_13_16,ip_14_15,p784,p785);
FA fa370(ip_15_14,ip_16_13,ip_17_12,p786,p787);
FA fa371(ip_18_11,ip_19_10,ip_20_9,p788,p789);
FA fa372(ip_21_8,ip_22_7,ip_23_6,p790,p791);
FA fa373(ip_24_5,ip_25_4,ip_26_3,p792,p793);
FA fa374(ip_27_2,ip_28_1,ip_29_0,p794,p795);
HA ha23(p777,p779,p796,p797);
FA fa375(p781,p783,p785,p798,p799);
FA fa376(p787,p789,p791,p800,p801);
FA fa377(p793,p795,p720,p802,p803);
FA fa378(p722,p724,p726,p804,p805);
FA fa379(p728,p730,p732,p806,p807);
FA fa380(p734,p736,p740,p808,p809);
FA fa381(p797,p738,p799,p810,p811);
FA fa382(p801,p803,p742,p812,p813);
FA fa383(p744,p805,p807,p814,p815);
FA fa384(p809,p746,p748,p816,p817);
FA fa385(p750,p752,p811,p818,p819);
FA fa386(p813,p754,p815,p820,p821);
FA fa387(p756,p758,p817,p822,p823);
FA fa388(p819,p760,p762,p824,p825);
FA fa389(p821,p764,p823,p826,p827);
FA fa390(p766,p825,p768,p828,p829);
FA fa391(p827,p770,p829,p830,p831);
FA fa392(p772,p831,p774,p832,p833);
FA fa393(ip_0_30,ip_1_29,ip_2_28,p834,p835);
FA fa394(ip_3_27,ip_4_26,ip_5_25,p836,p837);
FA fa395(ip_6_24,ip_7_23,ip_8_22,p838,p839);
FA fa396(ip_9_21,ip_10_20,ip_11_19,p840,p841);
FA fa397(ip_12_18,ip_13_17,ip_14_16,p842,p843);
FA fa398(ip_15_15,ip_16_14,ip_17_13,p844,p845);
FA fa399(ip_18_12,ip_19_11,ip_20_10,p846,p847);
FA fa400(ip_21_9,ip_22_8,ip_23_7,p848,p849);
FA fa401(ip_24_6,ip_25_5,ip_26_4,p850,p851);
FA fa402(ip_27_3,ip_28_2,ip_29_1,p852,p853);
FA fa403(ip_30_0,p835,p837,p854,p855);
FA fa404(p839,p841,p843,p856,p857);
FA fa405(p845,p847,p849,p858,p859);
FA fa406(p851,p853,p776,p860,p861);
FA fa407(p778,p780,p782,p862,p863);
FA fa408(p784,p786,p788,p864,p865);
FA fa409(p790,p792,p794,p866,p867);
FA fa410(p796,p855,p857,p868,p869);
FA fa411(p859,p861,p798,p870,p871);
FA fa412(p800,p802,p863,p872,p873);
FA fa413(p865,p867,p804,p874,p875);
FA fa414(p806,p808,p869,p876,p877);
FA fa415(p871,p810,p812,p878,p879);
FA fa416(p873,p875,p814,p880,p881);
FA fa417(p877,p816,p818,p882,p883);
FA fa418(p879,p881,p820,p884,p885);
FA fa419(p822,p883,p885,p886,p887);
FA fa420(p824,p826,p887,p888,p889);
FA fa421(p828,p889,p830,p890,p891);
FA fa422(ip_0_31,ip_1_30,ip_2_29,p892,p893);
FA fa423(ip_3_28,ip_4_27,ip_5_26,p894,p895);
FA fa424(ip_6_25,ip_7_24,ip_8_23,p896,p897);
FA fa425(ip_9_22,ip_10_21,ip_11_20,p898,p899);
FA fa426(ip_12_19,ip_13_18,ip_14_17,p900,p901);
FA fa427(ip_15_16,ip_16_15,ip_17_14,p902,p903);
FA fa428(ip_18_13,ip_19_12,ip_20_11,p904,p905);
FA fa429(ip_21_10,ip_22_9,ip_23_8,p906,p907);
FA fa430(ip_24_7,ip_25_6,ip_26_5,p908,p909);
FA fa431(ip_27_4,ip_28_3,ip_29_2,p910,p911);
FA fa432(ip_30_1,ip_31_0,p893,p912,p913);
FA fa433(p895,p897,p899,p914,p915);
FA fa434(p901,p903,p905,p916,p917);
FA fa435(p907,p909,p911,p918,p919);
FA fa436(p834,p836,p838,p920,p921);
FA fa437(p840,p842,p844,p922,p923);
FA fa438(p846,p848,p850,p924,p925);
FA fa439(p852,p913,p915,p926,p927);
FA fa440(p917,p919,p854,p928,p929);
FA fa441(p856,p858,p860,p930,p931);
FA fa442(p921,p923,p925,p932,p933);
FA fa443(p927,p862,p864,p934,p935);
FA fa444(p866,p929,p868,p936,p937);
FA fa445(p870,p931,p933,p938,p939);
FA fa446(p872,p874,p935,p940,p941);
FA fa447(p937,p876,p939,p942,p943);
FA fa448(p878,p880,p941,p944,p945);
FA fa449(p943,p882,p884,p946,p947);
HA ha24(p945,p886,p948,p949);
FA fa450(p947,p949,p888,p950,p951);
FA fa451(ip_1_31,ip_2_30,ip_3_29,p952,p953);
HA ha25(ip_4_28,ip_5_27,p954,p955);
FA fa452(ip_6_26,ip_7_25,ip_8_24,p956,p957);
FA fa453(ip_9_23,ip_10_22,ip_11_21,p958,p959);
FA fa454(ip_12_20,ip_13_19,ip_14_18,p960,p961);
FA fa455(ip_15_17,ip_16_16,ip_17_15,p962,p963);
FA fa456(ip_18_14,ip_19_13,ip_20_12,p964,p965);
FA fa457(ip_21_11,ip_22_10,ip_23_9,p966,p967);
FA fa458(ip_24_8,ip_25_7,ip_26_6,p968,p969);
FA fa459(ip_27_5,ip_28_4,ip_29_3,p970,p971);
FA fa460(ip_30_2,ip_31_1,p955,p972,p973);
FA fa461(p953,p957,p959,p974,p975);
FA fa462(p961,p963,p965,p976,p977);
FA fa463(p967,p969,p971,p978,p979);
FA fa464(p973,p892,p894,p980,p981);
FA fa465(p896,p898,p900,p982,p983);
HA ha26(p902,p904,p984,p985);
FA fa466(p906,p908,p910,p986,p987);
FA fa467(p912,p975,p977,p988,p989);
FA fa468(p979,p985,p914,p990,p991);
FA fa469(p916,p918,p981,p992,p993);
FA fa470(p983,p987,p920,p994,p995);
FA fa471(p922,p924,p926,p996,p997);
HA ha27(p989,p991,p998,p999);
FA fa472(p928,p993,p995,p1000,p1001);
FA fa473(p999,p930,p932,p1002,p1003);
FA fa474(p997,p1001,p934,p1004,p1005);
FA fa475(p936,p1003,p938,p1006,p1007);
FA fa476(p1005,p940,p1007,p1008,p1009);
FA fa477(p942,p1009,p944,p1010,p1011);
FA fa478(p1011,p946,p948,p1012,p1013);
FA fa479(ip_2_31,ip_3_30,ip_4_29,p1014,p1015);
FA fa480(ip_5_28,ip_6_27,ip_7_26,p1016,p1017);
FA fa481(ip_8_25,ip_9_24,ip_10_23,p1018,p1019);
HA ha28(ip_11_22,ip_12_21,p1020,p1021);
HA ha29(ip_13_20,ip_14_19,p1022,p1023);
HA ha30(ip_15_18,ip_16_17,p1024,p1025);
FA fa482(ip_17_16,ip_18_15,ip_19_14,p1026,p1027);
FA fa483(ip_20_13,ip_21_12,ip_22_11,p1028,p1029);
FA fa484(ip_23_10,ip_24_9,ip_25_8,p1030,p1031);
FA fa485(ip_26_7,ip_27_6,ip_28_5,p1032,p1033);
FA fa486(ip_29_4,ip_30_3,ip_31_2,p1034,p1035);
FA fa487(p1021,p1023,p1025,p1036,p1037);
HA ha31(p954,p1015,p1038,p1039);
FA fa488(p1017,p1019,p1027,p1040,p1041);
FA fa489(p1029,p1031,p1033,p1042,p1043);
FA fa490(p1035,p1037,p1039,p1044,p1045);
FA fa491(p952,p956,p958,p1046,p1047);
HA ha32(p960,p962,p1048,p1049);
FA fa492(p964,p966,p968,p1050,p1051);
FA fa493(p970,p972,p1041,p1052,p1053);
FA fa494(p1043,p1049,p984,p1054,p1055);
FA fa495(p1045,p1047,p1051,p1056,p1057);
FA fa496(p1053,p974,p976,p1058,p1059);
FA fa497(p978,p1055,p980,p1060,p1061);
FA fa498(p982,p986,p1057,p1062,p1063);
FA fa499(p1059,p988,p990,p1064,p1065);
FA fa500(p998,p1061,p1063,p1066,p1067);
HA ha33(p992,p994,p1068,p1069);
FA fa501(p1065,p1069,p996,p1070,p1071);
FA fa502(p1000,p1067,p1002,p1072,p1073);
FA fa503(p1071,p1004,p1073,p1074,p1075);
FA fa504(p1006,p1008,p1075,p1076,p1077);
FA fa505(p1010,p1077,p1012,p1078,p1079);
FA fa506(ip_3_31,ip_4_30,ip_5_29,p1080,p1081);
FA fa507(ip_6_28,ip_7_27,ip_8_26,p1082,p1083);
FA fa508(ip_9_25,ip_10_24,ip_11_23,p1084,p1085);
FA fa509(ip_12_22,ip_13_21,ip_14_20,p1086,p1087);
FA fa510(ip_15_19,ip_16_18,ip_17_17,p1088,p1089);
FA fa511(ip_18_16,ip_19_15,ip_20_14,p1090,p1091);
FA fa512(ip_21_13,ip_22_12,ip_23_11,p1092,p1093);
FA fa513(ip_24_10,ip_25_9,ip_26_8,p1094,p1095);
HA ha34(ip_27_7,ip_28_6,p1096,p1097);
FA fa514(ip_29_5,ip_30_4,ip_31_3,p1098,p1099);
FA fa515(p1020,p1022,p1024,p1100,p1101);
FA fa516(p1097,p1081,p1083,p1102,p1103);
FA fa517(p1085,p1087,p1089,p1104,p1105);
FA fa518(p1091,p1093,p1095,p1106,p1107);
FA fa519(p1099,p1014,p1016,p1108,p1109);
FA fa520(p1018,p1026,p1028,p1110,p1111);
FA fa521(p1030,p1032,p1034,p1112,p1113);
FA fa522(p1038,p1101,p1036,p1114,p1115);
FA fa523(p1048,p1103,p1105,p1116,p1117);
FA fa524(p1107,p1040,p1042,p1118,p1119);
FA fa525(p1109,p1111,p1113,p1120,p1121);
FA fa526(p1115,p1044,p1046,p1122,p1123);
FA fa527(p1050,p1052,p1117,p1124,p1125);
FA fa528(p1054,p1119,p1121,p1126,p1127);
FA fa529(p1056,p1058,p1123,p1128,p1129);
HA ha35(p1125,p1060,p1130,p1131);
HA ha36(p1062,p1068,p1132,p1133);
HA ha37(p1127,p1064,p1134,p1135);
FA fa530(p1129,p1131,p1133,p1136,p1137);
FA fa531(p1066,p1135,p1070,p1138,p1139);
FA fa532(p1137,p1072,p1139,p1140,p1141);
FA fa533(p1074,p1141,p1076,p1142,p1143);
FA fa534(ip_4_31,ip_5_30,ip_6_29,p1144,p1145);
FA fa535(ip_7_28,ip_8_27,ip_9_26,p1146,p1147);
FA fa536(ip_10_25,ip_11_24,ip_12_23,p1148,p1149);
FA fa537(ip_13_22,ip_14_21,ip_15_20,p1150,p1151);
FA fa538(ip_16_19,ip_17_18,ip_18_17,p1152,p1153);
FA fa539(ip_19_16,ip_20_15,ip_21_14,p1154,p1155);
FA fa540(ip_22_13,ip_23_12,ip_24_11,p1156,p1157);
FA fa541(ip_25_10,ip_26_9,ip_27_8,p1158,p1159);
HA ha38(ip_28_7,ip_29_6,p1160,p1161);
FA fa542(ip_30_5,ip_31_4,p1096,p1162,p1163);
FA fa543(p1161,p1145,p1147,p1164,p1165);
FA fa544(p1149,p1151,p1153,p1166,p1167);
FA fa545(p1155,p1157,p1159,p1168,p1169);
FA fa546(p1163,p1080,p1082,p1170,p1171);
FA fa547(p1084,p1086,p1088,p1172,p1173);
FA fa548(p1090,p1092,p1094,p1174,p1175);
FA fa549(p1098,p1100,p1165,p1176,p1177);
HA ha39(p1167,p1169,p1178,p1179);
FA fa550(p1102,p1104,p1106,p1180,p1181);
FA fa551(p1171,p1173,p1175,p1182,p1183);
FA fa552(p1179,p1108,p1110,p1184,p1185);
FA fa553(p1112,p1114,p1177,p1186,p1187);
FA fa554(p1116,p1181,p1183,p1188,p1189);
HA ha40(p1118,p1120,p1190,p1191);
FA fa555(p1185,p1187,p1122,p1192,p1193);
FA fa556(p1124,p1189,p1191,p1194,p1195);
HA ha41(p1126,p1130,p1196,p1197);
FA fa557(p1132,p1193,p1128,p1198,p1199);
FA fa558(p1134,p1195,p1197,p1200,p1201);
FA fa559(p1199,p1136,p1201,p1202,p1203);
FA fa560(p1138,p1203,p1140,p1204,p1205);
FA fa561(ip_5_31,ip_6_30,ip_7_29,p1206,p1207);
FA fa562(ip_8_28,ip_9_27,ip_10_26,p1208,p1209);
FA fa563(ip_11_25,ip_12_24,ip_13_23,p1210,p1211);
FA fa564(ip_14_22,ip_15_21,ip_16_20,p1212,p1213);
HA ha42(ip_17_19,ip_18_18,p1214,p1215);
FA fa565(ip_19_17,ip_20_16,ip_21_15,p1216,p1217);
FA fa566(ip_22_14,ip_23_13,ip_24_12,p1218,p1219);
FA fa567(ip_25_11,ip_26_10,ip_27_9,p1220,p1221);
FA fa568(ip_28_8,ip_29_7,ip_30_6,p1222,p1223);
FA fa569(ip_31_5,p1160,p1215,p1224,p1225);
HA ha43(p1207,p1209,p1226,p1227);
FA fa570(p1211,p1213,p1217,p1228,p1229);
FA fa571(p1219,p1221,p1223,p1230,p1231);
FA fa572(p1144,p1146,p1148,p1232,p1233);
FA fa573(p1150,p1152,p1154,p1234,p1235);
FA fa574(p1156,p1158,p1162,p1236,p1237);
FA fa575(p1225,p1227,p1229,p1238,p1239);
FA fa576(p1231,p1164,p1166,p1240,p1241);
FA fa577(p1168,p1178,p1233,p1242,p1243);
FA fa578(p1235,p1237,p1239,p1244,p1245);
FA fa579(p1170,p1172,p1174,p1246,p1247);
FA fa580(p1176,p1241,p1243,p1248,p1249);
FA fa581(p1245,p1180,p1182,p1250,p1251);
HA ha44(p1247,p1184,p1252,p1253);
FA fa582(p1186,p1190,p1249,p1254,p1255);
FA fa583(p1188,p1251,p1253,p1256,p1257);
FA fa584(p1192,p1196,p1255,p1258,p1259);
FA fa585(p1194,p1257,p1198,p1260,p1261);
FA fa586(p1259,p1200,p1261,p1262,p1263);
FA fa587(p1202,p1263,p1204,p1264,p1265);
FA fa588(ip_6_31,ip_7_30,ip_8_29,p1266,p1267);
FA fa589(ip_9_28,ip_10_27,ip_11_26,p1268,p1269);
FA fa590(ip_12_25,ip_13_24,ip_14_23,p1270,p1271);
FA fa591(ip_15_22,ip_16_21,ip_17_20,p1272,p1273);
FA fa592(ip_18_19,ip_19_18,ip_20_17,p1274,p1275);
FA fa593(ip_21_16,ip_22_15,ip_23_14,p1276,p1277);
FA fa594(ip_24_13,ip_25_12,ip_26_11,p1278,p1279);
FA fa595(ip_27_10,ip_28_9,ip_29_8,p1280,p1281);
FA fa596(ip_30_7,ip_31_6,p1214,p1282,p1283);
FA fa597(p1267,p1269,p1271,p1284,p1285);
FA fa598(p1273,p1275,p1277,p1286,p1287);
FA fa599(p1279,p1281,p1283,p1288,p1289);
FA fa600(p1206,p1208,p1210,p1290,p1291);
FA fa601(p1212,p1216,p1218,p1292,p1293);
FA fa602(p1220,p1222,p1226,p1294,p1295);
FA fa603(p1224,p1285,p1287,p1296,p1297);
FA fa604(p1289,p1228,p1230,p1298,p1299);
FA fa605(p1291,p1293,p1295,p1300,p1301);
FA fa606(p1232,p1234,p1236,p1302,p1303);
FA fa607(p1238,p1297,p1299,p1304,p1305);
FA fa608(p1301,p1240,p1242,p1306,p1307);
FA fa609(p1244,p1303,p1305,p1308,p1309);
FA fa610(p1246,p1248,p1252,p1310,p1311);
FA fa611(p1307,p1309,p1250,p1312,p1313);
HA ha45(p1254,p1311,p1314,p1315);
FA fa612(p1313,p1256,p1315,p1316,p1317);
FA fa613(p1258,p1260,p1317,p1318,p1319);
FA fa614(p1262,p1319,p1264,p1320,p1321);
FA fa615(ip_7_31,ip_8_30,ip_9_29,p1322,p1323);
FA fa616(ip_10_28,ip_11_27,ip_12_26,p1324,p1325);
FA fa617(ip_13_25,ip_14_24,ip_15_23,p1326,p1327);
FA fa618(ip_16_22,ip_17_21,ip_18_20,p1328,p1329);
FA fa619(ip_19_19,ip_20_18,ip_21_17,p1330,p1331);
FA fa620(ip_22_16,ip_23_15,ip_24_14,p1332,p1333);
FA fa621(ip_25_13,ip_26_12,ip_27_11,p1334,p1335);
FA fa622(ip_28_10,ip_29_9,ip_30_8,p1336,p1337);
FA fa623(ip_31_7,p1323,p1325,p1338,p1339);
FA fa624(p1327,p1329,p1331,p1340,p1341);
FA fa625(p1333,p1335,p1337,p1342,p1343);
FA fa626(p1266,p1268,p1270,p1344,p1345);
FA fa627(p1272,p1274,p1276,p1346,p1347);
FA fa628(p1278,p1280,p1282,p1348,p1349);
FA fa629(p1339,p1341,p1343,p1350,p1351);
FA fa630(p1284,p1286,p1288,p1352,p1353);
FA fa631(p1345,p1347,p1349,p1354,p1355);
FA fa632(p1290,p1292,p1294,p1356,p1357);
FA fa633(p1351,p1296,p1353,p1358,p1359);
FA fa634(p1355,p1298,p1300,p1360,p1361);
FA fa635(p1357,p1302,p1304,p1362,p1363);
FA fa636(p1359,p1361,p1306,p1364,p1365);
FA fa637(p1308,p1363,p1365,p1366,p1367);
FA fa638(p1310,p1312,p1314,p1368,p1369);
FA fa639(p1367,p1369,p1316,p1370,p1371);
FA fa640(p1371,p1318,p1320,p1372,p1373);
FA fa641(ip_8_31,ip_9_30,ip_10_29,p1374,p1375);
FA fa642(ip_11_28,ip_12_27,ip_13_26,p1376,p1377);
FA fa643(ip_14_25,ip_15_24,ip_16_23,p1378,p1379);
FA fa644(ip_17_22,ip_18_21,ip_19_20,p1380,p1381);
FA fa645(ip_20_19,ip_21_18,ip_22_17,p1382,p1383);
FA fa646(ip_23_16,ip_24_15,ip_25_14,p1384,p1385);
FA fa647(ip_26_13,ip_27_12,ip_28_11,p1386,p1387);
FA fa648(ip_29_10,ip_30_9,ip_31_8,p1388,p1389);
FA fa649(p1375,p1377,p1379,p1390,p1391);
FA fa650(p1381,p1383,p1385,p1392,p1393);
FA fa651(p1387,p1389,p1322,p1394,p1395);
FA fa652(p1324,p1326,p1328,p1396,p1397);
FA fa653(p1330,p1332,p1334,p1398,p1399);
FA fa654(p1336,p1391,p1393,p1400,p1401);
FA fa655(p1395,p1338,p1340,p1402,p1403);
FA fa656(p1342,p1397,p1399,p1404,p1405);
FA fa657(p1344,p1346,p1348,p1406,p1407);
FA fa658(p1401,p1350,p1403,p1408,p1409);
FA fa659(p1405,p1352,p1354,p1410,p1411);
FA fa660(p1407,p1356,p1409,p1412,p1413);
FA fa661(p1358,p1411,p1360,p1414,p1415);
FA fa662(p1413,p1362,p1415,p1416,p1417);
FA fa663(p1364,p1366,p1417,p1418,p1419);
FA fa664(p1368,p1419,p1370,p1420,p1421);
FA fa665(ip_9_31,ip_10_30,ip_11_29,p1422,p1423);
FA fa666(ip_12_28,ip_13_27,ip_14_26,p1424,p1425);
FA fa667(ip_15_25,ip_16_24,ip_17_23,p1426,p1427);
FA fa668(ip_18_22,ip_19_21,ip_20_20,p1428,p1429);
FA fa669(ip_21_19,ip_22_18,ip_23_17,p1430,p1431);
FA fa670(ip_24_16,ip_25_15,ip_26_14,p1432,p1433);
FA fa671(ip_27_13,ip_28_12,ip_29_11,p1434,p1435);
HA ha46(ip_30_10,ip_31_9,p1436,p1437);
FA fa672(p1437,p1423,p1425,p1438,p1439);
HA ha47(p1427,p1429,p1440,p1441);
FA fa673(p1431,p1433,p1435,p1442,p1443);
FA fa674(p1374,p1376,p1378,p1444,p1445);
FA fa675(p1380,p1382,p1384,p1446,p1447);
FA fa676(p1386,p1388,p1441,p1448,p1449);
FA fa677(p1439,p1443,p1390,p1450,p1451);
HA ha48(p1392,p1394,p1452,p1453);
FA fa678(p1445,p1447,p1449,p1454,p1455);
FA fa679(p1396,p1398,p1451,p1456,p1457);
FA fa680(p1453,p1400,p1455,p1458,p1459);
FA fa681(p1402,p1404,p1457,p1460,p1461);
FA fa682(p1406,p1459,p1408,p1462,p1463);
FA fa683(p1461,p1410,p1463,p1464,p1465);
FA fa684(p1412,p1414,p1465,p1466,p1467);
FA fa685(p1416,p1467,p1418,p1468,p1469);
HA ha49(ip_10_31,ip_11_30,p1470,p1471);
FA fa686(ip_12_29,ip_13_28,ip_14_27,p1472,p1473);
FA fa687(ip_15_26,ip_16_25,ip_17_24,p1474,p1475);
FA fa688(ip_18_23,ip_19_22,ip_20_21,p1476,p1477);
FA fa689(ip_21_20,ip_22_19,ip_23_18,p1478,p1479);
FA fa690(ip_24_17,ip_25_16,ip_26_15,p1480,p1481);
FA fa691(ip_27_14,ip_28_13,ip_29_12,p1482,p1483);
FA fa692(ip_30_11,ip_31_10,p1436,p1484,p1485);
FA fa693(p1471,p1473,p1475,p1486,p1487);
FA fa694(p1477,p1479,p1481,p1488,p1489);
FA fa695(p1483,p1485,p1422,p1490,p1491);
FA fa696(p1424,p1426,p1428,p1492,p1493);
FA fa697(p1430,p1432,p1434,p1494,p1495);
FA fa698(p1440,p1487,p1489,p1496,p1497);
FA fa699(p1491,p1438,p1442,p1498,p1499);
FA fa700(p1493,p1495,p1444,p1500,p1501);
FA fa701(p1446,p1448,p1452,p1502,p1503);
FA fa702(p1497,p1450,p1499,p1504,p1505);
FA fa703(p1501,p1454,p1503,p1506,p1507);
FA fa704(p1456,p1505,p1458,p1508,p1509);
FA fa705(p1507,p1460,p1509,p1510,p1511);
FA fa706(p1462,p1511,p1464,p1512,p1513);
FA fa707(p1513,p1466,p1468,p1514,p1515);
FA fa708(ip_11_31,ip_12_30,ip_13_29,p1516,p1517);
FA fa709(ip_14_28,ip_15_27,ip_16_26,p1518,p1519);
FA fa710(ip_17_25,ip_18_24,ip_19_23,p1520,p1521);
HA ha50(ip_20_22,ip_21_21,p1522,p1523);
FA fa711(ip_22_20,ip_23_19,ip_24_18,p1524,p1525);
FA fa712(ip_25_17,ip_26_16,ip_27_15,p1526,p1527);
FA fa713(ip_28_14,ip_29_13,ip_30_12,p1528,p1529);
FA fa714(ip_31_11,p1470,p1523,p1530,p1531);
FA fa715(p1517,p1519,p1521,p1532,p1533);
FA fa716(p1525,p1527,p1529,p1534,p1535);
FA fa717(p1472,p1474,p1476,p1536,p1537);
FA fa718(p1478,p1480,p1482,p1538,p1539);
HA ha51(p1484,p1531,p1540,p1541);
FA fa719(p1533,p1535,p1541,p1542,p1543);
FA fa720(p1486,p1488,p1490,p1544,p1545);
FA fa721(p1537,p1539,p1492,p1546,p1547);
FA fa722(p1494,p1543,p1496,p1548,p1549);
HA ha52(p1545,p1547,p1550,p1551);
FA fa723(p1498,p1500,p1549,p1552,p1553);
FA fa724(p1551,p1502,p1504,p1554,p1555);
FA fa725(p1553,p1506,p1555,p1556,p1557);
FA fa726(p1508,p1557,p1510,p1558,p1559);
FA fa727(p1559,p1512,p1514,p1560,p1561);
FA fa728(ip_12_31,ip_13_30,ip_14_29,p1562,p1563);
FA fa729(ip_15_28,ip_16_27,ip_17_26,p1564,p1565);
FA fa730(ip_18_25,ip_19_24,ip_20_23,p1566,p1567);
FA fa731(ip_21_22,ip_22_21,ip_23_20,p1568,p1569);
FA fa732(ip_24_19,ip_25_18,ip_26_17,p1570,p1571);
FA fa733(ip_27_16,ip_28_15,ip_29_14,p1572,p1573);
HA ha53(ip_30_13,ip_31_12,p1574,p1575);
FA fa734(p1522,p1575,p1563,p1576,p1577);
FA fa735(p1565,p1567,p1569,p1578,p1579);
FA fa736(p1571,p1573,p1516,p1580,p1581);
FA fa737(p1518,p1520,p1524,p1582,p1583);
FA fa738(p1526,p1528,p1577,p1584,p1585);
FA fa739(p1530,p1540,p1579,p1586,p1587);
FA fa740(p1581,p1532,p1534,p1588,p1589);
FA fa741(p1583,p1585,p1536,p1590,p1591);
FA fa742(p1538,p1587,p1542,p1592,p1593);
HA ha54(p1589,p1591,p1594,p1595);
FA fa743(p1544,p1546,p1550,p1596,p1597);
FA fa744(p1593,p1595,p1548,p1598,p1599);
FA fa745(p1597,p1599,p1552,p1600,p1601);
FA fa746(p1554,p1601,p1556,p1602,p1603);
HA ha55(p1603,p1558,p1604,p1605);
FA fa747(ip_13_31,ip_14_30,ip_15_29,p1606,p1607);
FA fa748(ip_16_28,ip_17_27,ip_18_26,p1608,p1609);
HA ha56(ip_19_25,ip_20_24,p1610,p1611);
FA fa749(ip_21_23,ip_22_22,ip_23_21,p1612,p1613);
FA fa750(ip_24_20,ip_25_19,ip_26_18,p1614,p1615);
HA ha57(ip_27_17,ip_28_16,p1616,p1617);
FA fa751(ip_29_15,ip_30_14,ip_31_13,p1618,p1619);
FA fa752(p1574,p1611,p1617,p1620,p1621);
HA ha58(p1607,p1609,p1622,p1623);
FA fa753(p1613,p1615,p1619,p1624,p1625);
FA fa754(p1562,p1564,p1566,p1626,p1627);
FA fa755(p1568,p1570,p1572,p1628,p1629);
FA fa756(p1621,p1623,p1576,p1630,p1631);
FA fa757(p1625,p1578,p1580,p1632,p1633);
FA fa758(p1627,p1629,p1631,p1634,p1635);
FA fa759(p1582,p1584,p1586,p1636,p1637);
FA fa760(p1633,p1635,p1588,p1638,p1639);
FA fa761(p1590,p1594,p1637,p1640,p1641);
FA fa762(p1592,p1639,p1641,p1642,p1643);
FA fa763(p1596,p1598,p1643,p1644,p1645);
FA fa764(p1600,p1645,p1602,p1646,p1647);
FA fa765(ip_14_31,ip_15_30,ip_16_29,p1648,p1649);
FA fa766(ip_17_28,ip_18_27,ip_19_26,p1650,p1651);
FA fa767(ip_20_25,ip_21_24,ip_22_23,p1652,p1653);
FA fa768(ip_23_22,ip_24_21,ip_25_20,p1654,p1655);
FA fa769(ip_26_19,ip_27_18,ip_28_17,p1656,p1657);
FA fa770(ip_29_16,ip_30_15,ip_31_14,p1658,p1659);
FA fa771(p1610,p1616,p1649,p1660,p1661);
FA fa772(p1651,p1653,p1655,p1662,p1663);
FA fa773(p1657,p1659,p1606,p1664,p1665);
FA fa774(p1608,p1612,p1614,p1666,p1667);
FA fa775(p1618,p1622,p1661,p1668,p1669);
FA fa776(p1620,p1663,p1665,p1670,p1671);
FA fa777(p1624,p1667,p1669,p1672,p1673);
FA fa778(p1626,p1628,p1630,p1674,p1675);
FA fa779(p1671,p1673,p1632,p1676,p1677);
FA fa780(p1634,p1675,p1636,p1678,p1679);
FA fa781(p1677,p1638,p1679,p1680,p1681);
FA fa782(p1640,p1642,p1681,p1682,p1683);
FA fa783(p1644,p1683,p1646,p1684,p1685);
FA fa784(ip_15_31,ip_16_30,ip_17_29,p1686,p1687);
FA fa785(ip_18_28,ip_19_27,ip_20_26,p1688,p1689);
FA fa786(ip_21_25,ip_22_24,ip_23_23,p1690,p1691);
FA fa787(ip_24_22,ip_25_21,ip_26_20,p1692,p1693);
FA fa788(ip_27_19,ip_28_18,ip_29_17,p1694,p1695);
FA fa789(ip_30_16,ip_31_15,p1687,p1696,p1697);
FA fa790(p1689,p1691,p1693,p1698,p1699);
FA fa791(p1695,p1648,p1650,p1700,p1701);
FA fa792(p1652,p1654,p1656,p1702,p1703);
FA fa793(p1658,p1697,p1660,p1704,p1705);
FA fa794(p1699,p1662,p1664,p1706,p1707);
FA fa795(p1701,p1703,p1705,p1708,p1709);
FA fa796(p1666,p1668,p1670,p1710,p1711);
FA fa797(p1707,p1709,p1672,p1712,p1713);
FA fa798(p1711,p1674,p1713,p1714,p1715);
FA fa799(p1676,p1678,p1715,p1716,p1717);
FA fa800(p1680,p1717,p1682,p1718,p1719);
FA fa801(ip_16_31,ip_17_30,ip_18_29,p1720,p1721);
FA fa802(ip_19_28,ip_20_27,ip_21_26,p1722,p1723);
FA fa803(ip_22_25,ip_23_24,ip_24_23,p1724,p1725);
HA ha59(ip_25_22,ip_26_21,p1726,p1727);
FA fa804(ip_27_20,ip_28_19,ip_29_18,p1728,p1729);
FA fa805(ip_30_17,ip_31_16,p1727,p1730,p1731);
FA fa806(p1721,p1723,p1725,p1732,p1733);
FA fa807(p1729,p1731,p1686,p1734,p1735);
FA fa808(p1688,p1690,p1692,p1736,p1737);
FA fa809(p1694,p1696,p1733,p1738,p1739);
FA fa810(p1735,p1698,p1737,p1740,p1741);
FA fa811(p1700,p1702,p1704,p1742,p1743);
FA fa812(p1739,p1741,p1706,p1744,p1745);
FA fa813(p1708,p1743,p1710,p1746,p1747);
HA ha60(p1745,p1712,p1748,p1749);
FA fa814(p1747,p1749,p1714,p1750,p1751);
FA fa815(p1751,p1716,p1718,p1752,p1753);
FA fa816(ip_17_31,ip_18_30,ip_19_29,p1754,p1755);
FA fa817(ip_20_28,ip_21_27,ip_22_26,p1756,p1757);
FA fa818(ip_23_25,ip_24_24,ip_25_23,p1758,p1759);
FA fa819(ip_26_22,ip_27_21,ip_28_20,p1760,p1761);
FA fa820(ip_29_19,ip_30_18,ip_31_17,p1762,p1763);
FA fa821(p1726,p1755,p1757,p1764,p1765);
FA fa822(p1759,p1761,p1763,p1766,p1767);
FA fa823(p1720,p1722,p1724,p1768,p1769);
FA fa824(p1728,p1730,p1765,p1770,p1771);
FA fa825(p1767,p1732,p1734,p1772,p1773);
FA fa826(p1769,p1771,p1736,p1774,p1775);
HA ha61(p1738,p1773,p1776,p1777);
FA fa827(p1775,p1740,p1777,p1778,p1779);
FA fa828(p1742,p1744,p1779,p1780,p1781);
FA fa829(p1746,p1748,p1781,p1782,p1783);
FA fa830(p1783,p1750,p1752,p1784,p1785);
FA fa831(ip_18_31,ip_19_30,ip_20_29,p1786,p1787);
FA fa832(ip_21_28,ip_22_27,ip_23_26,p1788,p1789);
FA fa833(ip_24_25,ip_25_24,ip_26_23,p1790,p1791);
FA fa834(ip_27_22,ip_28_21,ip_29_20,p1792,p1793);
HA ha62(ip_30_19,ip_31_18,p1794,p1795);
FA fa835(p1795,p1787,p1789,p1796,p1797);
HA ha63(p1791,p1793,p1798,p1799);
FA fa836(p1754,p1756,p1758,p1800,p1801);
FA fa837(p1760,p1762,p1799,p1802,p1803);
FA fa838(p1797,p1764,p1766,p1804,p1805);
FA fa839(p1801,p1803,p1768,p1806,p1807);
FA fa840(p1770,p1805,p1807,p1808,p1809);
FA fa841(p1772,p1774,p1776,p1810,p1811);
FA fa842(p1809,p1811,p1778,p1812,p1813);
FA fa843(p1813,p1780,p1782,p1814,p1815);
FA fa844(ip_19_31,ip_20_30,ip_21_29,p1816,p1817);
FA fa845(ip_22_28,ip_23_27,ip_24_26,p1818,p1819);
FA fa846(ip_25_25,ip_26_24,ip_27_23,p1820,p1821);
FA fa847(ip_28_22,ip_29_21,ip_30_20,p1822,p1823);
FA fa848(ip_31_19,p1794,p1817,p1824,p1825);
FA fa849(p1819,p1821,p1823,p1826,p1827);
FA fa850(p1786,p1788,p1790,p1828,p1829);
FA fa851(p1792,p1798,p1825,p1830,p1831);
FA fa852(p1827,p1796,p1829,p1832,p1833);
HA ha64(p1831,p1800,p1834,p1835);
FA fa853(p1802,p1833,p1835,p1836,p1837);
FA fa854(p1804,p1806,p1837,p1838,p1839);
FA fa855(p1808,p1839,p1810,p1840,p1841);
FA fa856(p1841,p1812,p1814,p1842,p1843);
HA ha65(ip_20_31,ip_21_30,p1844,p1845);
HA ha66(ip_22_29,ip_23_28,p1846,p1847);
FA fa857(ip_24_27,ip_25_26,ip_26_25,p1848,p1849);
FA fa858(ip_27_24,ip_28_23,ip_29_22,p1850,p1851);
FA fa859(ip_30_21,ip_31_20,p1845,p1852,p1853);
FA fa860(p1847,p1849,p1851,p1854,p1855);
FA fa861(p1853,p1816,p1818,p1856,p1857);
FA fa862(p1820,p1822,p1824,p1858,p1859);
FA fa863(p1855,p1826,p1857,p1860,p1861);
HA ha67(p1859,p1828,p1862,p1863);
FA fa864(p1830,p1834,p1861,p1864,p1865);
FA fa865(p1863,p1832,p1865,p1866,p1867);
FA fa866(p1836,p1867,p1838,p1868,p1869);
FA fa867(p1869,p1840,p1842,p1870,p1871);
FA fa868(ip_21_31,ip_22_30,ip_23_29,p1872,p1873);
FA fa869(ip_24_28,ip_25_27,ip_26_26,p1874,p1875);
FA fa870(ip_27_25,ip_28_24,ip_29_23,p1876,p1877);
FA fa871(ip_30_22,ip_31_21,p1844,p1878,p1879);
FA fa872(p1846,p1873,p1875,p1880,p1881);
HA ha68(p1877,p1879,p1882,p1883);
FA fa873(p1848,p1850,p1852,p1884,p1885);
FA fa874(p1883,p1881,p1854,p1886,p1887);
FA fa875(p1885,p1856,p1858,p1888,p1889);
FA fa876(p1887,p1862,p1860,p1890,p1891);
FA fa877(p1889,p1891,p1864,p1892,p1893);
FA fa878(p1866,p1893,p1868,p1894,p1895);
FA fa879(ip_22_31,ip_23_30,ip_24_29,p1896,p1897);
FA fa880(ip_25_28,ip_26_27,ip_27_26,p1898,p1899);
FA fa881(ip_28_25,ip_29_24,ip_30_23,p1900,p1901);
FA fa882(ip_31_22,p1897,p1899,p1902,p1903);
FA fa883(p1901,p1872,p1874,p1904,p1905);
FA fa884(p1876,p1878,p1882,p1906,p1907);
HA ha69(p1903,p1880,p1908,p1909);
FA fa885(p1905,p1907,p1884,p1910,p1911);
FA fa886(p1909,p1886,p1911,p1912,p1913);
HA ha70(p1888,p1913,p1914,p1915);
FA fa887(p1890,p1915,p1892,p1916,p1917);
FA fa888(ip_23_31,ip_24_30,ip_25_29,p1918,p1919);
FA fa889(ip_26_28,ip_27_27,ip_28_26,p1920,p1921);
FA fa890(ip_29_25,ip_30_24,ip_31_23,p1922,p1923);
FA fa891(p1919,p1921,p1923,p1924,p1925);
FA fa892(p1896,p1898,p1900,p1926,p1927);
FA fa893(p1925,p1902,p1927,p1928,p1929);
FA fa894(p1904,p1906,p1908,p1930,p1931);
FA fa895(p1929,p1910,p1931,p1932,p1933);
FA fa896(p1912,p1914,p1933,p1934,p1935);
FA fa897(ip_24_31,ip_25_30,ip_26_29,p1936,p1937);
HA ha71(ip_27_28,ip_28_27,p1938,p1939);
FA fa898(ip_29_26,ip_30_25,ip_31_24,p1940,p1941);
FA fa899(p1939,p1937,p1941,p1942,p1943);
FA fa900(p1918,p1920,p1922,p1944,p1945);
FA fa901(p1943,p1924,p1945,p1946,p1947);
FA fa902(p1926,p1947,p1928,p1948,p1949);
FA fa903(p1930,p1949,p1932,p1950,p1951);
FA fa904(ip_25_31,ip_26_30,ip_27_29,p1952,p1953);
FA fa905(ip_28_28,ip_29_27,ip_30_26,p1954,p1955);
FA fa906(ip_31_25,p1938,p1953,p1956,p1957);
FA fa907(p1955,p1936,p1940,p1958,p1959);
FA fa908(p1957,p1942,p1959,p1960,p1961);
FA fa909(p1944,p1961,p1946,p1962,p1963);
FA fa910(p1963,p1948,p1950,p1964,p1965);
FA fa911(ip_26_31,ip_27_30,ip_28_29,p1966,p1967);
FA fa912(ip_29_28,ip_30_27,ip_31_26,p1968,p1969);
FA fa913(p1967,p1969,p1952,p1970,p1971);
FA fa914(p1954,p1956,p1971,p1972,p1973);
FA fa915(p1958,p1973,p1960,p1974,p1975);
FA fa916(p1975,p1962,p1964,p1976,p1977);
FA fa917(ip_27_31,ip_28_30,ip_29_29,p1978,p1979);
FA fa918(ip_30_28,ip_31_27,p1979,p1980,p1981);
FA fa919(p1966,p1968,p1981,p1982,p1983);
HA ha72(p1970,p1983,p1984,p1985);
FA fa920(p1985,p1972,p1974,p1986,p1987);
HA ha73(ip_28_31,ip_29_30,p1988,p1989);
FA fa921(ip_30_29,ip_31_28,p1989,p1990,p1991);
FA fa922(p1991,p1978,p1980,p1992,p1993);
FA fa923(p1993,p1982,p1984,p1994,p1995);
FA fa924(ip_29_31,ip_30_30,ip_31_29,p1996,p1997);
FA fa925(p1988,p1997,p1990,p1998,p1999);
FA fa926(p1999,p1992,p1994,p2000,p2001);
FA fa927(ip_30_31,ip_31_30,p1996,p2002,p2003);
FA fa928(p2003,p1998,p2000,p2004,p2005);
HA ha74(ip_31_31,p2002,p2006,p2007);
wire [63:0] a,b;
wire [63:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p5;
assign b[3] = 1'b0;
assign a[4] = p11;
assign b[4] = 1'b0;
assign a[5] = p19;
assign b[5] = 1'b0;
assign a[6] = p29;
assign b[6] = 1'b0;
assign a[7] = p41;
assign b[7] = p28;
assign a[8] = p55;
assign b[8] = 1'b0;
assign a[9] = p71;
assign b[9] = 1'b0;
assign a[10] = p89;
assign b[10] = p70;
assign a[11] = p109;
assign b[11] = p88;
assign a[12] = p108;
assign b[12] = p131;
assign a[13] = p155;
assign b[13] = p130;
assign a[14] = p181;
assign b[14] = p154;
assign a[15] = p211;
assign b[15] = p180;
assign a[16] = p243;
assign b[16] = 1'b0;
assign a[17] = p277;
assign b[17] = 1'b0;
assign a[18] = p311;
assign b[18] = p276;
assign a[19] = p349;
assign b[19] = 1'b0;
assign a[20] = p389;
assign b[20] = 1'b0;
assign a[21] = p429;
assign b[21] = p388;
assign a[22] = p471;
assign b[22] = 1'b0;
assign a[23] = p515;
assign b[23] = 1'b0;
assign a[24] = p563;
assign b[24] = p514;
assign a[25] = p613;
assign b[25] = 1'b0;
assign a[26] = p665;
assign b[26] = p612;
assign a[27] = p719;
assign b[27] = p664;
assign a[28] = p775;
assign b[28] = 1'b0;
assign a[29] = p833;
assign b[29] = 1'b0;
assign a[30] = p891;
assign b[30] = p832;
assign a[31] = p951;
assign b[31] = p890;
assign a[32] = p1013;
assign b[32] = p950;
assign a[33] = p1079;
assign b[33] = 1'b0;
assign a[34] = p1143;
assign b[34] = p1078;
assign a[35] = p1205;
assign b[35] = p1142;
assign a[36] = p1265;
assign b[36] = 1'b0;
assign a[37] = p1321;
assign b[37] = 1'b0;
assign a[38] = p1373;
assign b[38] = 1'b0;
assign a[39] = p1421;
assign b[39] = p1372;
assign a[40] = p1469;
assign b[40] = p1420;
assign a[41] = p1515;
assign b[41] = 1'b0;
assign a[42] = p1561;
assign b[42] = 1'b0;
assign a[43] = p1605;
assign b[43] = p1560;
assign a[44] = p1604;
assign b[44] = p1647;
assign a[45] = p1685;
assign b[45] = 1'b0;
assign a[46] = p1719;
assign b[46] = p1684;
assign a[47] = p1753;
assign b[47] = 1'b0;
assign a[48] = p1785;
assign b[48] = 1'b0;
assign a[49] = p1815;
assign b[49] = p1784;
assign a[50] = p1843;
assign b[50] = 1'b0;
assign a[51] = p1871;
assign b[51] = 1'b0;
assign a[52] = p1895;
assign b[52] = p1870;
assign a[53] = p1917;
assign b[53] = p1894;
assign a[54] = p1935;
assign b[54] = p1916;
assign a[55] = p1951;
assign b[55] = p1934;
assign a[56] = p1965;
assign b[56] = 1'b0;
assign a[57] = p1977;
assign b[57] = 1'b0;
assign a[58] = p1987;
assign b[58] = p1976;
assign a[59] = p1995;
assign b[59] = p1986;
assign a[60] = p2001;
assign b[60] = 1'b0;
assign a[61] = p2005;
assign b[61] = 1'b0;
assign a[62] = p2007;
assign b[62] = p2004;
assign a[63] = p2006;
assign b[63] = 1'b0;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[63] = s[63];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
assign o[31] = s[31];
assign o[32] = s[32];
assign o[33] = s[33];
assign o[34] = s[34];
assign o[35] = s[35];
assign o[36] = s[36];
assign o[37] = s[37];
assign o[38] = s[38];
assign o[39] = s[39];
assign o[40] = s[40];
assign o[41] = s[41];
assign o[42] = s[42];
assign o[43] = s[43];
assign o[44] = s[44];
assign o[45] = s[45];
assign o[46] = s[46];
assign o[47] = s[47];
assign o[48] = s[48];
assign o[49] = s[49];
assign o[50] = s[50];
assign o[51] = s[51];
assign o[52] = s[52];
assign o[53] = s[53];
assign o[54] = s[54];
assign o[55] = s[55];
assign o[56] = s[56];
assign o[57] = s[57];
assign o[58] = s[58];
assign o[59] = s[59];
assign o[60] = s[60];
assign o[61] = s[61];
assign o[62] = s[62];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [63:0] a,b;
output [63:0] s;
assign s = a+b;
endmodule
