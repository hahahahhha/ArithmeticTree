// 1 2 2 2 2 2 1 2 1 2 2 2 2 1 2 2 1 2 1 2 2 1 2 2 1 2 2 2 2 1 2 3 

module main(x,y,o);
input [15:0] x,y;
output [31:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_1_0,x[1],y[0]);
and and17(ip_1_1,x[1],y[1]);
and and18(ip_1_2,x[1],y[2]);
and and19(ip_1_3,x[1],y[3]);
and and20(ip_1_4,x[1],y[4]);
and and21(ip_1_5,x[1],y[5]);
and and22(ip_1_6,x[1],y[6]);
and and23(ip_1_7,x[1],y[7]);
and and24(ip_1_8,x[1],y[8]);
and and25(ip_1_9,x[1],y[9]);
and and26(ip_1_10,x[1],y[10]);
and and27(ip_1_11,x[1],y[11]);
and and28(ip_1_12,x[1],y[12]);
and and29(ip_1_13,x[1],y[13]);
and and30(ip_1_14,x[1],y[14]);
and and31(ip_1_15,x[1],y[15]);
and and32(ip_2_0,x[2],y[0]);
and and33(ip_2_1,x[2],y[1]);
and and34(ip_2_2,x[2],y[2]);
and and35(ip_2_3,x[2],y[3]);
and and36(ip_2_4,x[2],y[4]);
and and37(ip_2_5,x[2],y[5]);
and and38(ip_2_6,x[2],y[6]);
and and39(ip_2_7,x[2],y[7]);
and and40(ip_2_8,x[2],y[8]);
and and41(ip_2_9,x[2],y[9]);
and and42(ip_2_10,x[2],y[10]);
and and43(ip_2_11,x[2],y[11]);
and and44(ip_2_12,x[2],y[12]);
and and45(ip_2_13,x[2],y[13]);
and and46(ip_2_14,x[2],y[14]);
and and47(ip_2_15,x[2],y[15]);
and and48(ip_3_0,x[3],y[0]);
and and49(ip_3_1,x[3],y[1]);
and and50(ip_3_2,x[3],y[2]);
and and51(ip_3_3,x[3],y[3]);
and and52(ip_3_4,x[3],y[4]);
and and53(ip_3_5,x[3],y[5]);
and and54(ip_3_6,x[3],y[6]);
and and55(ip_3_7,x[3],y[7]);
and and56(ip_3_8,x[3],y[8]);
and and57(ip_3_9,x[3],y[9]);
and and58(ip_3_10,x[3],y[10]);
and and59(ip_3_11,x[3],y[11]);
and and60(ip_3_12,x[3],y[12]);
and and61(ip_3_13,x[3],y[13]);
and and62(ip_3_14,x[3],y[14]);
and and63(ip_3_15,x[3],y[15]);
and and64(ip_4_0,x[4],y[0]);
and and65(ip_4_1,x[4],y[1]);
and and66(ip_4_2,x[4],y[2]);
and and67(ip_4_3,x[4],y[3]);
and and68(ip_4_4,x[4],y[4]);
and and69(ip_4_5,x[4],y[5]);
and and70(ip_4_6,x[4],y[6]);
and and71(ip_4_7,x[4],y[7]);
and and72(ip_4_8,x[4],y[8]);
and and73(ip_4_9,x[4],y[9]);
and and74(ip_4_10,x[4],y[10]);
and and75(ip_4_11,x[4],y[11]);
and and76(ip_4_12,x[4],y[12]);
and and77(ip_4_13,x[4],y[13]);
and and78(ip_4_14,x[4],y[14]);
and and79(ip_4_15,x[4],y[15]);
and and80(ip_5_0,x[5],y[0]);
and and81(ip_5_1,x[5],y[1]);
and and82(ip_5_2,x[5],y[2]);
and and83(ip_5_3,x[5],y[3]);
and and84(ip_5_4,x[5],y[4]);
and and85(ip_5_5,x[5],y[5]);
and and86(ip_5_6,x[5],y[6]);
and and87(ip_5_7,x[5],y[7]);
and and88(ip_5_8,x[5],y[8]);
and and89(ip_5_9,x[5],y[9]);
and and90(ip_5_10,x[5],y[10]);
and and91(ip_5_11,x[5],y[11]);
and and92(ip_5_12,x[5],y[12]);
and and93(ip_5_13,x[5],y[13]);
and and94(ip_5_14,x[5],y[14]);
and and95(ip_5_15,x[5],y[15]);
and and96(ip_6_0,x[6],y[0]);
and and97(ip_6_1,x[6],y[1]);
and and98(ip_6_2,x[6],y[2]);
and and99(ip_6_3,x[6],y[3]);
and and100(ip_6_4,x[6],y[4]);
and and101(ip_6_5,x[6],y[5]);
and and102(ip_6_6,x[6],y[6]);
and and103(ip_6_7,x[6],y[7]);
and and104(ip_6_8,x[6],y[8]);
and and105(ip_6_9,x[6],y[9]);
and and106(ip_6_10,x[6],y[10]);
and and107(ip_6_11,x[6],y[11]);
and and108(ip_6_12,x[6],y[12]);
and and109(ip_6_13,x[6],y[13]);
and and110(ip_6_14,x[6],y[14]);
and and111(ip_6_15,x[6],y[15]);
and and112(ip_7_0,x[7],y[0]);
and and113(ip_7_1,x[7],y[1]);
and and114(ip_7_2,x[7],y[2]);
and and115(ip_7_3,x[7],y[3]);
and and116(ip_7_4,x[7],y[4]);
and and117(ip_7_5,x[7],y[5]);
and and118(ip_7_6,x[7],y[6]);
and and119(ip_7_7,x[7],y[7]);
and and120(ip_7_8,x[7],y[8]);
and and121(ip_7_9,x[7],y[9]);
and and122(ip_7_10,x[7],y[10]);
and and123(ip_7_11,x[7],y[11]);
and and124(ip_7_12,x[7],y[12]);
and and125(ip_7_13,x[7],y[13]);
and and126(ip_7_14,x[7],y[14]);
and and127(ip_7_15,x[7],y[15]);
and and128(ip_8_0,x[8],y[0]);
and and129(ip_8_1,x[8],y[1]);
and and130(ip_8_2,x[8],y[2]);
and and131(ip_8_3,x[8],y[3]);
and and132(ip_8_4,x[8],y[4]);
and and133(ip_8_5,x[8],y[5]);
and and134(ip_8_6,x[8],y[6]);
and and135(ip_8_7,x[8],y[7]);
and and136(ip_8_8,x[8],y[8]);
and and137(ip_8_9,x[8],y[9]);
and and138(ip_8_10,x[8],y[10]);
and and139(ip_8_11,x[8],y[11]);
and and140(ip_8_12,x[8],y[12]);
and and141(ip_8_13,x[8],y[13]);
and and142(ip_8_14,x[8],y[14]);
and and143(ip_8_15,x[8],y[15]);
and and144(ip_9_0,x[9],y[0]);
and and145(ip_9_1,x[9],y[1]);
and and146(ip_9_2,x[9],y[2]);
and and147(ip_9_3,x[9],y[3]);
and and148(ip_9_4,x[9],y[4]);
and and149(ip_9_5,x[9],y[5]);
and and150(ip_9_6,x[9],y[6]);
and and151(ip_9_7,x[9],y[7]);
and and152(ip_9_8,x[9],y[8]);
and and153(ip_9_9,x[9],y[9]);
and and154(ip_9_10,x[9],y[10]);
and and155(ip_9_11,x[9],y[11]);
and and156(ip_9_12,x[9],y[12]);
and and157(ip_9_13,x[9],y[13]);
and and158(ip_9_14,x[9],y[14]);
and and159(ip_9_15,x[9],y[15]);
and and160(ip_10_0,x[10],y[0]);
and and161(ip_10_1,x[10],y[1]);
and and162(ip_10_2,x[10],y[2]);
and and163(ip_10_3,x[10],y[3]);
and and164(ip_10_4,x[10],y[4]);
and and165(ip_10_5,x[10],y[5]);
and and166(ip_10_6,x[10],y[6]);
and and167(ip_10_7,x[10],y[7]);
and and168(ip_10_8,x[10],y[8]);
and and169(ip_10_9,x[10],y[9]);
and and170(ip_10_10,x[10],y[10]);
and and171(ip_10_11,x[10],y[11]);
and and172(ip_10_12,x[10],y[12]);
and and173(ip_10_13,x[10],y[13]);
and and174(ip_10_14,x[10],y[14]);
and and175(ip_10_15,x[10],y[15]);
and and176(ip_11_0,x[11],y[0]);
and and177(ip_11_1,x[11],y[1]);
and and178(ip_11_2,x[11],y[2]);
and and179(ip_11_3,x[11],y[3]);
and and180(ip_11_4,x[11],y[4]);
and and181(ip_11_5,x[11],y[5]);
and and182(ip_11_6,x[11],y[6]);
and and183(ip_11_7,x[11],y[7]);
and and184(ip_11_8,x[11],y[8]);
and and185(ip_11_9,x[11],y[9]);
and and186(ip_11_10,x[11],y[10]);
and and187(ip_11_11,x[11],y[11]);
and and188(ip_11_12,x[11],y[12]);
and and189(ip_11_13,x[11],y[13]);
and and190(ip_11_14,x[11],y[14]);
and and191(ip_11_15,x[11],y[15]);
and and192(ip_12_0,x[12],y[0]);
and and193(ip_12_1,x[12],y[1]);
and and194(ip_12_2,x[12],y[2]);
and and195(ip_12_3,x[12],y[3]);
and and196(ip_12_4,x[12],y[4]);
and and197(ip_12_5,x[12],y[5]);
and and198(ip_12_6,x[12],y[6]);
and and199(ip_12_7,x[12],y[7]);
and and200(ip_12_8,x[12],y[8]);
and and201(ip_12_9,x[12],y[9]);
and and202(ip_12_10,x[12],y[10]);
and and203(ip_12_11,x[12],y[11]);
and and204(ip_12_12,x[12],y[12]);
and and205(ip_12_13,x[12],y[13]);
and and206(ip_12_14,x[12],y[14]);
and and207(ip_12_15,x[12],y[15]);
and and208(ip_13_0,x[13],y[0]);
and and209(ip_13_1,x[13],y[1]);
and and210(ip_13_2,x[13],y[2]);
and and211(ip_13_3,x[13],y[3]);
and and212(ip_13_4,x[13],y[4]);
and and213(ip_13_5,x[13],y[5]);
and and214(ip_13_6,x[13],y[6]);
and and215(ip_13_7,x[13],y[7]);
and and216(ip_13_8,x[13],y[8]);
and and217(ip_13_9,x[13],y[9]);
and and218(ip_13_10,x[13],y[10]);
and and219(ip_13_11,x[13],y[11]);
and and220(ip_13_12,x[13],y[12]);
and and221(ip_13_13,x[13],y[13]);
and and222(ip_13_14,x[13],y[14]);
and and223(ip_13_15,x[13],y[15]);
and and224(ip_14_0,x[14],y[0]);
and and225(ip_14_1,x[14],y[1]);
and and226(ip_14_2,x[14],y[2]);
and and227(ip_14_3,x[14],y[3]);
and and228(ip_14_4,x[14],y[4]);
and and229(ip_14_5,x[14],y[5]);
and and230(ip_14_6,x[14],y[6]);
and and231(ip_14_7,x[14],y[7]);
and and232(ip_14_8,x[14],y[8]);
and and233(ip_14_9,x[14],y[9]);
and and234(ip_14_10,x[14],y[10]);
and and235(ip_14_11,x[14],y[11]);
and and236(ip_14_12,x[14],y[12]);
and and237(ip_14_13,x[14],y[13]);
and and238(ip_14_14,x[14],y[14]);
and and239(ip_14_15,x[14],y[15]);
and and240(ip_15_0,x[15],y[0]);
and and241(ip_15_1,x[15],y[1]);
and and242(ip_15_2,x[15],y[2]);
and and243(ip_15_3,x[15],y[3]);
and and244(ip_15_4,x[15],y[4]);
and and245(ip_15_5,x[15],y[5]);
and and246(ip_15_6,x[15],y[6]);
and and247(ip_15_7,x[15],y[7]);
and and248(ip_15_8,x[15],y[8]);
and and249(ip_15_9,x[15],y[9]);
and and250(ip_15_10,x[15],y[10]);
and and251(ip_15_11,x[15],y[11]);
and and252(ip_15_12,x[15],y[12]);
and and253(ip_15_13,x[15],y[13]);
and and254(ip_15_14,x[15],y[14]);
and and255(ip_15_15,x[15],y[15]);
HA ha0(ip_0_2,ip_1_1,p0,p1);
FA fa0(ip_0_3,ip_1_2,ip_2_1,p2,p3);
HA ha1(ip_3_0,p0,p4,p5);
FA fa1(ip_0_4,ip_1_3,ip_2_2,p6,p7);
FA fa2(ip_3_1,ip_4_0,p4,p8,p9);
HA ha2(p7,p2,p10,p11);
FA fa3(ip_0_5,ip_1_4,ip_2_3,p12,p13);
HA ha3(ip_3_2,ip_4_1,p14,p15);
FA fa4(ip_5_0,p15,p13,p16,p17);
HA ha4(p17,p6,p18,p19);
HA ha5(p10,p19,p20,p21);
FA fa5(ip_0_6,ip_1_5,ip_2_4,p22,p23);
FA fa6(ip_3_3,ip_4_2,ip_5_1,p24,p25);
HA ha6(ip_6_0,p14,p26,p27);
FA fa7(p23,p25,p27,p28,p29);
FA fa8(p12,p16,p18,p30,p31);
FA fa9(p29,p20,p31,p32,p33);
FA fa10(ip_0_7,ip_1_6,ip_2_5,p34,p35);
HA ha7(ip_3_4,ip_4_3,p36,p37);
FA fa11(ip_5_2,ip_6_1,ip_7_0,p38,p39);
FA fa12(p37,p26,p35,p40,p41);
FA fa13(p39,p22,p24,p42,p43);
FA fa14(p41,p28,p43,p44,p45);
HA ha8(p30,p45,p46,p47);
HA ha9(ip_0_8,ip_1_7,p48,p49);
HA ha10(ip_2_6,ip_3_5,p50,p51);
FA fa15(ip_4_4,ip_5_3,ip_6_2,p52,p53);
HA ha11(ip_7_1,ip_8_0,p54,p55);
FA fa16(p36,p49,p51,p56,p57);
FA fa17(p55,p53,p34,p58,p59);
FA fa18(p38,p57,p59,p60,p61);
HA ha12(p40,p61,p62,p63);
HA ha13(p42,p63,p64,p65);
FA fa19(p65,p44,p46,p66,p67);
FA fa20(ip_0_9,ip_1_8,ip_2_7,p68,p69);
HA ha14(ip_3_6,ip_4_5,p70,p71);
FA fa21(ip_5_4,ip_6_3,ip_7_2,p72,p73);
FA fa22(ip_8_1,ip_9_0,p48,p74,p75);
FA fa23(p50,p54,p71,p76,p77);
FA fa24(p69,p73,p75,p78,p79);
HA ha15(p52,p77,p80,p81);
FA fa25(p56,p79,p81,p82,p83);
HA ha16(p58,p60,p84,p85);
HA ha17(p62,p83,p86,p87);
FA fa26(p64,p85,p87,p88,p89);
FA fa27(ip_0_10,ip_1_9,ip_2_8,p90,p91);
HA ha18(ip_3_7,ip_4_6,p92,p93);
HA ha19(ip_5_5,ip_6_4,p94,p95);
HA ha20(ip_7_3,ip_8_2,p96,p97);
HA ha21(ip_9_1,ip_10_0,p98,p99);
HA ha22(p70,p93,p100,p101);
HA ha23(p95,p97,p102,p103);
FA fa28(p99,p101,p103,p104,p105);
HA ha24(p91,p68,p106,p107);
HA ha25(p72,p74,p108,p109);
HA ha26(p105,p107,p110,p111);
HA ha27(p109,p76,p112,p113);
FA fa29(p80,p111,p113,p114,p115);
FA fa30(p78,p115,p82,p116,p117);
HA ha28(p84,p86,p118,p119);
HA ha29(p119,p117,p120,p121);
FA fa31(ip_0_11,ip_1_10,ip_2_9,p122,p123);
FA fa32(ip_3_8,ip_4_7,ip_5_6,p124,p125);
FA fa33(ip_6_5,ip_7_4,ip_8_3,p126,p127);
HA ha30(ip_9_2,ip_10_1,p128,p129);
HA ha31(ip_11_0,p129,p130,p131);
HA ha32(p92,p94,p132,p133);
HA ha33(p96,p98,p134,p135);
HA ha34(p100,p102,p136,p137);
FA fa34(p123,p125,p127,p138,p139);
HA ha35(p131,p133,p140,p141);
HA ha36(p135,p137,p142,p143);
HA ha37(p141,p90,p144,p145);
FA fa35(p106,p108,p139,p146,p147);
FA fa36(p143,p145,p104,p148,p149);
FA fa37(p110,p112,p147,p150,p151);
HA ha38(p149,p151,p152,p153);
HA ha39(p114,p118,p154,p155);
FA fa38(p153,p155,p116,p156,p157);
HA ha40(ip_0_12,ip_1_11,p158,p159);
HA ha41(ip_2_10,ip_3_9,p160,p161);
HA ha42(ip_4_8,ip_5_7,p162,p163);
HA ha43(ip_6_6,ip_7_5,p164,p165);
HA ha44(ip_8_4,ip_9_3,p166,p167);
HA ha45(ip_10_2,ip_11_1,p168,p169);
HA ha46(ip_12_0,p128,p170,p171);
FA fa39(p159,p161,p163,p172,p173);
HA ha47(p165,p167,p174,p175);
HA ha48(p169,p130,p176,p177);
HA ha49(p132,p134,p178,p179);
FA fa40(p171,p175,p122,p180,p181);
HA ha50(p124,p126,p182,p183);
FA fa41(p136,p140,p173,p184,p185);
FA fa42(p177,p179,p142,p186,p187);
FA fa43(p144,p181,p183,p188,p189);
FA fa44(p138,p185,p187,p190,p191);
HA ha51(p189,p146,p192,p193);
FA fa45(p148,p191,p150,p194,p195);
HA ha52(p152,p193,p196,p197);
FA fa46(p154,p195,p197,p198,p199);
FA fa47(ip_0_13,ip_1_12,ip_2_11,p200,p201);
FA fa48(ip_3_10,ip_4_9,ip_5_8,p202,p203);
FA fa49(ip_6_7,ip_7_6,ip_8_5,p204,p205);
HA ha53(ip_9_4,ip_10_3,p206,p207);
FA fa50(ip_11_2,ip_12_1,ip_13_0,p208,p209);
FA fa51(p158,p160,p162,p210,p211);
FA fa52(p164,p166,p168,p212,p213);
FA fa53(p207,p170,p174,p214,p215);
FA fa54(p201,p203,p205,p216,p217);
FA fa55(p209,p176,p178,p218,p219);
FA fa56(p211,p213,p172,p220,p221);
HA ha54(p182,p215,p222,p223);
FA fa57(p217,p180,p219,p224,p225);
FA fa58(p221,p223,p184,p226,p227);
HA ha55(p186,p188,p228,p229);
FA fa59(p225,p227,p190,p230,p231);
HA ha56(p192,p229,p232,p233);
FA fa60(p196,p231,p233,p234,p235);
FA fa61(p194,p235,p198,p236,p237);
HA ha57(ip_0_14,ip_1_13,p238,p239);
HA ha58(ip_2_12,ip_3_11,p240,p241);
HA ha59(ip_4_10,ip_5_9,p242,p243);
HA ha60(ip_6_8,ip_7_7,p244,p245);
HA ha61(ip_8_6,ip_9_5,p246,p247);
FA fa62(ip_10_4,ip_11_3,ip_12_2,p248,p249);
FA fa63(ip_13_1,ip_14_0,p206,p250,p251);
FA fa64(p239,p241,p243,p252,p253);
HA ha62(p245,p247,p254,p255);
FA fa65(p249,p251,p255,p256,p257);
FA fa66(p200,p202,p204,p258,p259);
FA fa67(p208,p253,p210,p260,p261);
HA ha63(p212,p257,p262,p263);
HA ha64(p214,p216,p264,p265);
FA fa68(p222,p259,p261,p266,p267);
FA fa69(p263,p218,p220,p268,p269);
HA ha65(p265,p267,p270,p271);
FA fa70(p224,p226,p228,p272,p273);
FA fa71(p269,p271,p232,p274,p275);
FA fa72(p230,p273,p275,p276,p277);
HA ha66(p234,p277,p278,p279);
FA fa73(ip_0_15,ip_1_14,ip_2_13,p280,p281);
FA fa74(ip_3_12,ip_4_11,ip_5_10,p282,p283);
FA fa75(ip_6_9,ip_7_8,ip_8_7,p284,p285);
FA fa76(ip_9_6,ip_10_5,ip_11_4,p286,p287);
FA fa77(ip_12_3,ip_13_2,ip_14_1,p288,p289);
FA fa78(ip_15_0,p238,p240,p290,p291);
HA ha67(p242,p244,p292,p293);
HA ha68(p246,p254,p294,p295);
FA fa79(p281,p283,p285,p296,p297);
FA fa80(p287,p289,p293,p298,p299);
FA fa81(p248,p250,p291,p300,p301);
HA ha69(p295,p252,p302,p303);
HA ha70(p297,p299,p304,p305);
HA ha71(p256,p262,p306,p307);
FA fa82(p301,p303,p305,p308,p309);
HA ha72(p258,p260,p310,p311);
HA ha73(p264,p307,p312,p313);
HA ha74(p309,p311,p314,p315);
HA ha75(p313,p266,p316,p317);
HA ha76(p270,p315,p318,p319);
FA fa83(p268,p317,p319,p320,p321);
FA fa84(p272,p274,p321,p322,p323);
HA ha77(p276,p278,p324,p325);
FA fa85(ip_1_15,ip_2_14,ip_3_13,p326,p327);
FA fa86(ip_4_12,ip_5_11,ip_6_10,p328,p329);
HA ha78(ip_7_9,ip_8_8,p330,p331);
FA fa87(ip_9_7,ip_10_6,ip_11_5,p332,p333);
HA ha79(ip_12_4,ip_13_3,p334,p335);
HA ha80(ip_14_2,ip_15_1,p336,p337);
HA ha81(p331,p335,p338,p339);
FA fa88(p337,p292,p327,p340,p341);
FA fa89(p329,p333,p339,p342,p343);
FA fa90(p280,p282,p284,p344,p345);
FA fa91(p286,p288,p294,p346,p347);
HA ha82(p290,p341,p348,p349);
HA ha83(p343,p296,p350,p351);
FA fa92(p298,p302,p304,p352,p353);
HA ha84(p345,p347,p354,p355);
FA fa93(p349,p300,p306,p356,p357);
HA ha85(p351,p355,p358,p359);
HA ha86(p310,p312,p360,p361);
FA fa94(p353,p359,p308,p362,p363);
HA ha87(p314,p357,p364,p365);
FA fa95(p361,p316,p318,p366,p367);
FA fa96(p363,p365,p367,p368,p369);
HA ha88(p320,p369,p370,p371);
FA fa97(p371,p322,p324,p372,p373);
HA ha89(ip_2_15,ip_3_14,p374,p375);
FA fa98(ip_4_13,ip_5_12,ip_6_11,p376,p377);
FA fa99(ip_7_10,ip_8_9,ip_9_8,p378,p379);
HA ha90(ip_10_7,ip_11_6,p380,p381);
HA ha91(ip_12_5,ip_13_4,p382,p383);
HA ha92(ip_14_3,ip_15_2,p384,p385);
FA fa100(p330,p334,p336,p386,p387);
FA fa101(p375,p381,p383,p388,p389);
FA fa102(p385,p338,p377,p390,p391);
FA fa103(p379,p326,p328,p392,p393);
FA fa104(p332,p387,p389,p394,p395);
HA ha93(p391,p340,p396,p397);
FA fa105(p342,p348,p393,p398,p399);
FA fa106(p395,p344,p346,p400,p401);
HA ha94(p350,p354,p402,p403);
FA fa107(p397,p358,p399,p404,p405);
FA fa108(p403,p352,p360,p406,p407);
FA fa109(p401,p356,p364,p408,p409);
FA fa110(p405,p362,p407,p410,p411);
FA fa111(p409,p366,p411,p412,p413);
FA fa112(p368,p370,p413,p414,p415);
FA fa113(ip_3_15,ip_4_14,ip_5_13,p416,p417);
FA fa114(ip_6_12,ip_7_11,ip_8_10,p418,p419);
FA fa115(ip_9_9,ip_10_8,ip_11_7,p420,p421);
FA fa116(ip_12_6,ip_13_5,ip_14_4,p422,p423);
HA ha95(ip_15_3,p374,p424,p425);
HA ha96(p380,p382,p426,p427);
FA fa117(p384,p417,p419,p428,p429);
FA fa118(p421,p423,p425,p430,p431);
FA fa119(p427,p376,p378,p432,p433);
FA fa120(p386,p388,p429,p434,p435);
FA fa121(p431,p390,p433,p436,p437);
HA ha97(p392,p394,p438,p439);
FA fa122(p396,p435,p402,p440,p441);
FA fa123(p437,p439,p398,p442,p443);
FA fa124(p441,p400,p443,p444,p445);
HA ha98(p404,p406,p446,p447);
FA fa125(p445,p408,p447,p448,p449);
HA ha99(p410,p449,p450,p451);
FA fa126(p412,p451,p414,p452,p453);
FA fa127(ip_4_15,ip_5_14,ip_6_13,p454,p455);
HA ha100(ip_7_12,ip_8_11,p456,p457);
FA fa128(ip_9_10,ip_10_9,ip_11_8,p458,p459);
HA ha101(ip_12_7,ip_13_6,p460,p461);
HA ha102(ip_14_5,ip_15_4,p462,p463);
FA fa129(p457,p461,p463,p464,p465);
HA ha103(p424,p426,p466,p467);
FA fa130(p455,p459,p416,p468,p469);
FA fa131(p418,p420,p422,p470,p471);
FA fa132(p465,p467,p469,p472,p473);
FA fa133(p428,p430,p471,p474,p475);
HA ha104(p473,p432,p476,p477);
FA fa134(p434,p438,p475,p478,p479);
FA fa135(p477,p436,p440,p480,p481);
FA fa136(p479,p442,p481,p482,p483);
FA fa137(p444,p446,p483,p484,p485);
FA fa138(p485,p448,p450,p486,p487);
HA ha105(ip_5_15,ip_6_14,p488,p489);
FA fa139(ip_7_13,ip_8_12,ip_9_11,p490,p491);
HA ha106(ip_10_10,ip_11_9,p492,p493);
HA ha107(ip_12_8,ip_13_7,p494,p495);
FA fa140(ip_14_6,ip_15_5,p456,p496,p497);
FA fa141(p460,p462,p489,p498,p499);
HA ha108(p493,p495,p500,p501);
HA ha109(p491,p497,p502,p503);
FA fa142(p501,p454,p458,p504,p505);
FA fa143(p466,p499,p503,p506,p507);
FA fa144(p464,p468,p505,p508,p509);
HA ha110(p507,p470,p510,p511);
FA fa145(p472,p476,p509,p512,p513);
HA ha111(p511,p474,p514,p515);
HA ha112(p513,p515,p516,p517);
HA ha113(p478,p517,p518,p519);
HA ha114(p480,p519,p520,p521);
FA fa146(p521,p482,p484,p522,p523);
HA ha115(ip_6_15,ip_7_14,p524,p525);
FA fa147(ip_8_13,ip_9_12,ip_10_11,p526,p527);
HA ha116(ip_11_10,ip_12_9,p528,p529);
HA ha117(ip_13_8,ip_14_7,p530,p531);
FA fa148(ip_15_6,p488,p492,p532,p533);
HA ha118(p494,p525,p534,p535);
HA ha119(p529,p531,p536,p537);
HA ha120(p500,p527,p538,p539);
HA ha121(p535,p537,p540,p541);
HA ha122(p490,p496,p542,p543);
FA fa149(p502,p533,p539,p544,p545);
HA ha123(p541,p498,p546,p547);
FA fa150(p543,p545,p547,p548,p549);
FA fa151(p504,p506,p510,p550,p551);
HA ha124(p549,p508,p552,p553);
FA fa152(p551,p514,p553,p554,p555);
FA fa153(p512,p516,p518,p556,p557);
HA ha125(p555,p520,p558,p559);
FA fa154(p557,p559,p522,p560,p561);
FA fa155(ip_7_15,ip_8_14,ip_9_13,p562,p563);
FA fa156(ip_10_12,ip_11_11,ip_12_10,p564,p565);
HA ha126(ip_13_9,ip_14_8,p566,p567);
HA ha127(ip_15_7,p524,p568,p569);
HA ha128(p528,p530,p570,p571);
HA ha129(p567,p534,p572,p573);
FA fa157(p536,p563,p565,p574,p575);
HA ha130(p569,p571,p576,p577);
HA ha131(p526,p538,p578,p579);
HA ha132(p540,p573,p580,p581);
FA fa158(p577,p532,p542,p582,p583);
HA ha133(p575,p579,p584,p585);
HA ha134(p581,p546,p586,p587);
FA fa159(p585,p544,p583,p588,p589);
FA fa160(p587,p548,p589,p590,p591);
HA ha135(p550,p552,p592,p593);
FA fa161(p591,p593,p554,p594,p595);
FA fa162(p556,p558,p595,p596,p597);
HA ha136(ip_8_15,ip_9_14,p598,p599);
FA fa163(ip_10_13,ip_11_12,ip_12_11,p600,p601);
FA fa164(ip_13_10,ip_14_9,ip_15_8,p602,p603);
FA fa165(p566,p599,p568,p604,p605);
HA ha137(p570,p601,p606,p607);
FA fa166(p603,p562,p564,p608,p609);
HA ha138(p572,p576,p610,p611);
HA ha139(p605,p607,p612,p613);
HA ha140(p578,p580,p614,p615);
HA ha141(p611,p613,p616,p617);
HA ha142(p574,p584,p618,p619);
FA fa167(p609,p615,p617,p620,p621);
FA fa168(p586,p619,p582,p622,p623);
FA fa169(p621,p623,p588,p624,p625);
FA fa170(p592,p625,p590,p626,p627);
HA ha143(p627,p594,p628,p629);
FA fa171(ip_9_15,ip_10_14,ip_11_13,p630,p631);
FA fa172(ip_12_12,ip_13_11,ip_14_10,p632,p633);
HA ha144(ip_15_9,p598,p634,p635);
FA fa173(p631,p633,p635,p636,p637);
FA fa174(p600,p602,p606,p638,p639);
FA fa175(p604,p610,p612,p640,p641);
FA fa176(p637,p614,p616,p642,p643);
FA fa177(p639,p608,p618,p644,p645);
FA fa178(p641,p643,p620,p646,p647);
HA ha145(p645,p622,p648,p649);
FA fa179(p647,p649,p624,p650,p651);
FA fa180(p651,p626,p628,p652,p653);
FA fa181(ip_10_15,ip_11_14,ip_12_13,p654,p655);
HA ha146(ip_13_12,ip_14_11,p656,p657);
FA fa182(ip_15_10,p657,p634,p658,p659);
FA fa183(p655,p630,p632,p660,p661);
HA ha147(p659,p636,p662,p663);
HA ha148(p661,p638,p664,p665);
FA fa184(p663,p640,p665,p666,p667);
FA fa185(p642,p644,p667,p668,p669);
FA fa186(p646,p648,p669,p670,p671);
HA ha149(p671,p650,p672,p673);
FA fa187(ip_11_15,ip_12_14,ip_13_13,p674,p675);
FA fa188(ip_14_12,ip_15_11,p656,p676,p677);
HA ha150(p675,p677,p678,p679);
FA fa189(p654,p679,p658,p680,p681);
HA ha151(p681,p660,p682,p683);
HA ha152(p662,p664,p684,p685);
FA fa190(p683,p685,p666,p686,p687);
FA fa191(p687,p668,p670,p688,p689);
FA fa192(ip_12_15,ip_13_14,ip_14_13,p690,p691);
FA fa193(ip_15_12,p691,p674,p692,p693);
HA ha153(p676,p678,p694,p695);
FA fa194(p693,p695,p680,p696,p697);
HA ha154(p682,p697,p698,p699);
FA fa195(p684,p699,p686,p700,p701);
FA fa196(ip_13_15,ip_14_14,ip_15_13,p702,p703);
HA ha155(p703,p690,p704,p705);
FA fa197(p694,p705,p692,p706,p707);
HA ha156(p707,p696,p708,p709);
HA ha157(p698,p709,p710,p711);
HA ha158(ip_14_15,ip_15_14,p712,p713);
HA ha159(p713,p702,p714,p715);
FA fa198(p704,p715,p706,p716,p717);
FA fa199(p717,p708,p710,p718,p719);
HA ha160(ip_15_15,p712,p720,p721);
HA ha161(p721,p714,p722,p723);
HA ha162(p723,p716,p724,p725);
wire [31:0] a,b;
wire [31:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = ip_2_0;
assign b[2] = p1;
assign a[3] = p3;
assign b[3] = p5;
assign a[4] = p9;
assign b[4] = p11;
assign a[5] = p8;
assign b[5] = p21;
assign a[6] = p33;
assign b[6] = 1'b0;
assign a[7] = p32;
assign b[7] = p47;
assign a[8] = p67;
assign b[8] = 1'b0;
assign a[9] = p89;
assign b[9] = p66;
assign a[10] = p121;
assign b[10] = p88;
assign a[11] = p120;
assign b[11] = p157;
assign a[12] = p199;
assign b[12] = p156;
assign a[13] = p237;
assign b[13] = 1'b0;
assign a[14] = p279;
assign b[14] = p236;
assign a[15] = p323;
assign b[15] = p325;
assign a[16] = p373;
assign b[16] = 1'b0;
assign a[17] = p415;
assign b[17] = p372;
assign a[18] = p453;
assign b[18] = 1'b0;
assign a[19] = p487;
assign b[19] = p452;
assign a[20] = p523;
assign b[20] = p486;
assign a[21] = p561;
assign b[21] = 1'b0;
assign a[22] = p597;
assign b[22] = p560;
assign a[23] = p629;
assign b[23] = p596;
assign a[24] = p653;
assign b[24] = 1'b0;
assign a[25] = p673;
assign b[25] = p652;
assign a[26] = p672;
assign b[26] = p689;
assign a[27] = p701;
assign b[27] = p688;
assign a[28] = p711;
assign b[28] = p700;
assign a[29] = p719;
assign b[29] = 1'b0;
assign a[30] = p725;
assign b[30] = p718;
assign a[31] = p720;
assign b[31] = p722;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[31] = s[31] & p724;
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [31:0] a,b;
output [31:0] s;
assign s = a+b;
endmodule
