// 1 2 1 1 2 2 2 2 1 2 2 2 2 2 2 2 1 2 2 2 2 1 1 2 2 2 1 1 1 2 2 1 

module main(x,y,o);
input [15:0] x,y;
output [31:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_1_0,x[1],y[0]);
and and17(ip_1_1,x[1],y[1]);
and and18(ip_1_2,x[1],y[2]);
and and19(ip_1_3,x[1],y[3]);
and and20(ip_1_4,x[1],y[4]);
and and21(ip_1_5,x[1],y[5]);
and and22(ip_1_6,x[1],y[6]);
and and23(ip_1_7,x[1],y[7]);
and and24(ip_1_8,x[1],y[8]);
and and25(ip_1_9,x[1],y[9]);
and and26(ip_1_10,x[1],y[10]);
and and27(ip_1_11,x[1],y[11]);
and and28(ip_1_12,x[1],y[12]);
and and29(ip_1_13,x[1],y[13]);
and and30(ip_1_14,x[1],y[14]);
and and31(ip_1_15,x[1],y[15]);
and and32(ip_2_0,x[2],y[0]);
and and33(ip_2_1,x[2],y[1]);
and and34(ip_2_2,x[2],y[2]);
and and35(ip_2_3,x[2],y[3]);
and and36(ip_2_4,x[2],y[4]);
and and37(ip_2_5,x[2],y[5]);
and and38(ip_2_6,x[2],y[6]);
and and39(ip_2_7,x[2],y[7]);
and and40(ip_2_8,x[2],y[8]);
and and41(ip_2_9,x[2],y[9]);
and and42(ip_2_10,x[2],y[10]);
and and43(ip_2_11,x[2],y[11]);
and and44(ip_2_12,x[2],y[12]);
and and45(ip_2_13,x[2],y[13]);
and and46(ip_2_14,x[2],y[14]);
and and47(ip_2_15,x[2],y[15]);
and and48(ip_3_0,x[3],y[0]);
and and49(ip_3_1,x[3],y[1]);
and and50(ip_3_2,x[3],y[2]);
and and51(ip_3_3,x[3],y[3]);
and and52(ip_3_4,x[3],y[4]);
and and53(ip_3_5,x[3],y[5]);
and and54(ip_3_6,x[3],y[6]);
and and55(ip_3_7,x[3],y[7]);
and and56(ip_3_8,x[3],y[8]);
and and57(ip_3_9,x[3],y[9]);
and and58(ip_3_10,x[3],y[10]);
and and59(ip_3_11,x[3],y[11]);
and and60(ip_3_12,x[3],y[12]);
and and61(ip_3_13,x[3],y[13]);
and and62(ip_3_14,x[3],y[14]);
and and63(ip_3_15,x[3],y[15]);
and and64(ip_4_0,x[4],y[0]);
and and65(ip_4_1,x[4],y[1]);
and and66(ip_4_2,x[4],y[2]);
and and67(ip_4_3,x[4],y[3]);
and and68(ip_4_4,x[4],y[4]);
and and69(ip_4_5,x[4],y[5]);
and and70(ip_4_6,x[4],y[6]);
and and71(ip_4_7,x[4],y[7]);
and and72(ip_4_8,x[4],y[8]);
and and73(ip_4_9,x[4],y[9]);
and and74(ip_4_10,x[4],y[10]);
and and75(ip_4_11,x[4],y[11]);
and and76(ip_4_12,x[4],y[12]);
and and77(ip_4_13,x[4],y[13]);
and and78(ip_4_14,x[4],y[14]);
and and79(ip_4_15,x[4],y[15]);
and and80(ip_5_0,x[5],y[0]);
and and81(ip_5_1,x[5],y[1]);
and and82(ip_5_2,x[5],y[2]);
and and83(ip_5_3,x[5],y[3]);
and and84(ip_5_4,x[5],y[4]);
and and85(ip_5_5,x[5],y[5]);
and and86(ip_5_6,x[5],y[6]);
and and87(ip_5_7,x[5],y[7]);
and and88(ip_5_8,x[5],y[8]);
and and89(ip_5_9,x[5],y[9]);
and and90(ip_5_10,x[5],y[10]);
and and91(ip_5_11,x[5],y[11]);
and and92(ip_5_12,x[5],y[12]);
and and93(ip_5_13,x[5],y[13]);
and and94(ip_5_14,x[5],y[14]);
and and95(ip_5_15,x[5],y[15]);
and and96(ip_6_0,x[6],y[0]);
and and97(ip_6_1,x[6],y[1]);
and and98(ip_6_2,x[6],y[2]);
and and99(ip_6_3,x[6],y[3]);
and and100(ip_6_4,x[6],y[4]);
and and101(ip_6_5,x[6],y[5]);
and and102(ip_6_6,x[6],y[6]);
and and103(ip_6_7,x[6],y[7]);
and and104(ip_6_8,x[6],y[8]);
and and105(ip_6_9,x[6],y[9]);
and and106(ip_6_10,x[6],y[10]);
and and107(ip_6_11,x[6],y[11]);
and and108(ip_6_12,x[6],y[12]);
and and109(ip_6_13,x[6],y[13]);
and and110(ip_6_14,x[6],y[14]);
and and111(ip_6_15,x[6],y[15]);
and and112(ip_7_0,x[7],y[0]);
and and113(ip_7_1,x[7],y[1]);
and and114(ip_7_2,x[7],y[2]);
and and115(ip_7_3,x[7],y[3]);
and and116(ip_7_4,x[7],y[4]);
and and117(ip_7_5,x[7],y[5]);
and and118(ip_7_6,x[7],y[6]);
and and119(ip_7_7,x[7],y[7]);
and and120(ip_7_8,x[7],y[8]);
and and121(ip_7_9,x[7],y[9]);
and and122(ip_7_10,x[7],y[10]);
and and123(ip_7_11,x[7],y[11]);
and and124(ip_7_12,x[7],y[12]);
and and125(ip_7_13,x[7],y[13]);
and and126(ip_7_14,x[7],y[14]);
and and127(ip_7_15,x[7],y[15]);
and and128(ip_8_0,x[8],y[0]);
and and129(ip_8_1,x[8],y[1]);
and and130(ip_8_2,x[8],y[2]);
and and131(ip_8_3,x[8],y[3]);
and and132(ip_8_4,x[8],y[4]);
and and133(ip_8_5,x[8],y[5]);
and and134(ip_8_6,x[8],y[6]);
and and135(ip_8_7,x[8],y[7]);
and and136(ip_8_8,x[8],y[8]);
and and137(ip_8_9,x[8],y[9]);
and and138(ip_8_10,x[8],y[10]);
and and139(ip_8_11,x[8],y[11]);
and and140(ip_8_12,x[8],y[12]);
and and141(ip_8_13,x[8],y[13]);
and and142(ip_8_14,x[8],y[14]);
and and143(ip_8_15,x[8],y[15]);
and and144(ip_9_0,x[9],y[0]);
and and145(ip_9_1,x[9],y[1]);
and and146(ip_9_2,x[9],y[2]);
and and147(ip_9_3,x[9],y[3]);
and and148(ip_9_4,x[9],y[4]);
and and149(ip_9_5,x[9],y[5]);
and and150(ip_9_6,x[9],y[6]);
and and151(ip_9_7,x[9],y[7]);
and and152(ip_9_8,x[9],y[8]);
and and153(ip_9_9,x[9],y[9]);
and and154(ip_9_10,x[9],y[10]);
and and155(ip_9_11,x[9],y[11]);
and and156(ip_9_12,x[9],y[12]);
and and157(ip_9_13,x[9],y[13]);
and and158(ip_9_14,x[9],y[14]);
and and159(ip_9_15,x[9],y[15]);
and and160(ip_10_0,x[10],y[0]);
and and161(ip_10_1,x[10],y[1]);
and and162(ip_10_2,x[10],y[2]);
and and163(ip_10_3,x[10],y[3]);
and and164(ip_10_4,x[10],y[4]);
and and165(ip_10_5,x[10],y[5]);
and and166(ip_10_6,x[10],y[6]);
and and167(ip_10_7,x[10],y[7]);
and and168(ip_10_8,x[10],y[8]);
and and169(ip_10_9,x[10],y[9]);
and and170(ip_10_10,x[10],y[10]);
and and171(ip_10_11,x[10],y[11]);
and and172(ip_10_12,x[10],y[12]);
and and173(ip_10_13,x[10],y[13]);
and and174(ip_10_14,x[10],y[14]);
and and175(ip_10_15,x[10],y[15]);
and and176(ip_11_0,x[11],y[0]);
and and177(ip_11_1,x[11],y[1]);
and and178(ip_11_2,x[11],y[2]);
and and179(ip_11_3,x[11],y[3]);
and and180(ip_11_4,x[11],y[4]);
and and181(ip_11_5,x[11],y[5]);
and and182(ip_11_6,x[11],y[6]);
and and183(ip_11_7,x[11],y[7]);
and and184(ip_11_8,x[11],y[8]);
and and185(ip_11_9,x[11],y[9]);
and and186(ip_11_10,x[11],y[10]);
and and187(ip_11_11,x[11],y[11]);
and and188(ip_11_12,x[11],y[12]);
and and189(ip_11_13,x[11],y[13]);
and and190(ip_11_14,x[11],y[14]);
and and191(ip_11_15,x[11],y[15]);
and and192(ip_12_0,x[12],y[0]);
and and193(ip_12_1,x[12],y[1]);
and and194(ip_12_2,x[12],y[2]);
and and195(ip_12_3,x[12],y[3]);
and and196(ip_12_4,x[12],y[4]);
and and197(ip_12_5,x[12],y[5]);
and and198(ip_12_6,x[12],y[6]);
and and199(ip_12_7,x[12],y[7]);
and and200(ip_12_8,x[12],y[8]);
and and201(ip_12_9,x[12],y[9]);
and and202(ip_12_10,x[12],y[10]);
and and203(ip_12_11,x[12],y[11]);
and and204(ip_12_12,x[12],y[12]);
and and205(ip_12_13,x[12],y[13]);
and and206(ip_12_14,x[12],y[14]);
and and207(ip_12_15,x[12],y[15]);
and and208(ip_13_0,x[13],y[0]);
and and209(ip_13_1,x[13],y[1]);
and and210(ip_13_2,x[13],y[2]);
and and211(ip_13_3,x[13],y[3]);
and and212(ip_13_4,x[13],y[4]);
and and213(ip_13_5,x[13],y[5]);
and and214(ip_13_6,x[13],y[6]);
and and215(ip_13_7,x[13],y[7]);
and and216(ip_13_8,x[13],y[8]);
and and217(ip_13_9,x[13],y[9]);
and and218(ip_13_10,x[13],y[10]);
and and219(ip_13_11,x[13],y[11]);
and and220(ip_13_12,x[13],y[12]);
and and221(ip_13_13,x[13],y[13]);
and and222(ip_13_14,x[13],y[14]);
and and223(ip_13_15,x[13],y[15]);
and and224(ip_14_0,x[14],y[0]);
and and225(ip_14_1,x[14],y[1]);
and and226(ip_14_2,x[14],y[2]);
and and227(ip_14_3,x[14],y[3]);
and and228(ip_14_4,x[14],y[4]);
and and229(ip_14_5,x[14],y[5]);
and and230(ip_14_6,x[14],y[6]);
and and231(ip_14_7,x[14],y[7]);
and and232(ip_14_8,x[14],y[8]);
and and233(ip_14_9,x[14],y[9]);
and and234(ip_14_10,x[14],y[10]);
and and235(ip_14_11,x[14],y[11]);
and and236(ip_14_12,x[14],y[12]);
and and237(ip_14_13,x[14],y[13]);
and and238(ip_14_14,x[14],y[14]);
and and239(ip_14_15,x[14],y[15]);
and and240(ip_15_0,x[15],y[0]);
and and241(ip_15_1,x[15],y[1]);
and and242(ip_15_2,x[15],y[2]);
and and243(ip_15_3,x[15],y[3]);
and and244(ip_15_4,x[15],y[4]);
and and245(ip_15_5,x[15],y[5]);
and and246(ip_15_6,x[15],y[6]);
and and247(ip_15_7,x[15],y[7]);
and and248(ip_15_8,x[15],y[8]);
and and249(ip_15_9,x[15],y[9]);
and and250(ip_15_10,x[15],y[10]);
and and251(ip_15_11,x[15],y[11]);
and and252(ip_15_12,x[15],y[12]);
and and253(ip_15_13,x[15],y[13]);
and and254(ip_15_14,x[15],y[14]);
and and255(ip_15_15,x[15],y[15]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
FA fa2(ip_3_0,p3,p0,p4,p5);
HA ha0(ip_0_4,ip_1_3,p6,p7);
FA fa3(ip_2_2,ip_3_1,ip_4_0,p8,p9);
FA fa4(p7,p9,p2,p10,p11);
FA fa5(ip_0_5,ip_1_4,ip_2_3,p12,p13);
HA ha1(ip_3_2,ip_4_1,p14,p15);
FA fa6(ip_5_0,p15,p6,p16,p17);
FA fa7(p13,p17,p8,p18,p19);
HA ha2(ip_0_6,ip_1_5,p20,p21);
FA fa8(ip_2_4,ip_3_3,ip_4_2,p22,p23);
FA fa9(ip_5_1,ip_6_0,p14,p24,p25);
FA fa10(p21,p23,p25,p26,p27);
FA fa11(p12,p16,p27,p28,p29);
FA fa12(ip_0_7,ip_1_6,ip_2_5,p30,p31);
FA fa13(ip_3_4,ip_4_3,ip_5_2,p32,p33);
HA ha3(ip_6_1,ip_7_0,p34,p35);
HA ha4(p20,p35,p36,p37);
HA ha5(p31,p33,p38,p39);
FA fa14(p37,p22,p24,p40,p41);
FA fa15(p39,p26,p41,p42,p43);
FA fa16(ip_0_8,ip_1_7,ip_2_6,p44,p45);
FA fa17(ip_3_5,ip_4_4,ip_5_3,p46,p47);
FA fa18(ip_6_2,ip_7_1,ip_8_0,p48,p49);
FA fa19(p34,p36,p45,p50,p51);
HA ha6(p47,p49,p52,p53);
FA fa20(p30,p32,p38,p54,p55);
FA fa21(p53,p51,p55,p56,p57);
FA fa22(p40,p57,p42,p58,p59);
FA fa23(ip_0_9,ip_1_8,ip_2_7,p60,p61);
HA ha7(ip_3_6,ip_4_5,p62,p63);
FA fa24(ip_5_4,ip_6_3,ip_7_2,p64,p65);
FA fa25(ip_8_1,ip_9_0,p63,p66,p67);
FA fa26(p61,p65,p67,p68,p69);
HA ha8(p44,p46,p70,p71);
HA ha9(p48,p52,p72,p73);
FA fa27(p69,p71,p73,p74,p75);
FA fa28(p50,p54,p75,p76,p77);
HA ha10(p56,p77,p78,p79);
HA ha11(ip_0_10,ip_1_9,p80,p81);
FA fa29(ip_2_8,ip_3_7,ip_4_6,p82,p83);
FA fa30(ip_5_5,ip_6_4,ip_7_3,p84,p85);
HA ha12(ip_8_2,ip_9_1,p86,p87);
FA fa31(ip_10_0,p62,p81,p88,p89);
FA fa32(p87,p83,p85,p90,p91);
HA ha13(p60,p64,p92,p93);
FA fa33(p66,p89,p70,p94,p95);
FA fa34(p72,p91,p93,p96,p97);
FA fa35(p68,p95,p97,p98,p99);
HA ha14(p74,p99,p100,p101);
HA ha15(p101,p76,p102,p103);
FA fa36(ip_0_11,ip_1_10,ip_2_9,p104,p105);
FA fa37(ip_3_8,ip_4_7,ip_5_6,p106,p107);
HA ha16(ip_6_5,ip_7_4,p108,p109);
FA fa38(ip_8_3,ip_9_2,ip_10_1,p110,p111);
HA ha17(ip_11_0,p109,p112,p113);
HA ha18(p80,p86,p114,p115);
FA fa39(p105,p107,p111,p116,p117);
FA fa40(p113,p115,p82,p118,p119);
FA fa41(p84,p117,p119,p120,p121);
HA ha19(p88,p92,p122,p123);
FA fa42(p123,p90,p121,p124,p125);
HA ha20(p94,p125,p126,p127);
HA ha21(p96,p100,p128,p129);
HA ha22(p127,p98,p130,p131);
HA ha23(p129,p131,p132,p133);
FA fa43(ip_0_12,ip_1_11,ip_2_10,p134,p135);
FA fa44(ip_3_9,ip_4_8,ip_5_7,p136,p137);
FA fa45(ip_6_6,ip_7_5,ip_8_4,p138,p139);
FA fa46(ip_9_3,ip_10_2,ip_11_1,p140,p141);
HA ha24(ip_12_0,p108,p142,p143);
HA ha25(p112,p114,p144,p145);
FA fa47(p135,p137,p139,p146,p147);
HA ha26(p141,p143,p148,p149);
FA fa48(p104,p106,p110,p150,p151);
FA fa49(p145,p149,p147,p152,p153);
HA ha27(p116,p118,p154,p155);
FA fa50(p122,p151,p153,p156,p157);
FA fa51(p155,p120,p157,p158,p159);
FA fa52(p124,p126,p128,p160,p161);
FA fa53(p130,p159,p132,p162,p163);
HA ha28(ip_0_13,ip_1_12,p164,p165);
HA ha29(ip_2_11,ip_3_10,p166,p167);
HA ha30(ip_4_9,ip_5_8,p168,p169);
HA ha31(ip_6_7,ip_7_6,p170,p171);
FA fa54(ip_8_5,ip_9_4,ip_10_3,p172,p173);
HA ha32(ip_11_2,ip_12_1,p174,p175);
FA fa55(ip_13_0,p165,p167,p176,p177);
FA fa56(p169,p171,p175,p178,p179);
HA ha33(p142,p173,p180,p181);
HA ha34(p134,p136,p182,p183);
HA ha35(p138,p140,p184,p185);
FA fa57(p144,p148,p177,p186,p187);
HA ha36(p179,p181,p188,p189);
HA ha37(p183,p185,p190,p191);
FA fa58(p189,p146,p187,p192,p193);
HA ha38(p191,p150,p194,p195);
FA fa59(p152,p154,p193,p196,p197);
HA ha39(p195,p156,p198,p199);
FA fa60(p197,p199,p158,p200,p201);
HA ha40(p160,p201,p202,p203);
HA ha41(ip_0_14,ip_1_13,p204,p205);
HA ha42(ip_2_12,ip_3_11,p206,p207);
FA fa61(ip_4_10,ip_5_9,ip_6_8,p208,p209);
HA ha43(ip_7_7,ip_8_6,p210,p211);
HA ha44(ip_9_5,ip_10_4,p212,p213);
HA ha45(ip_11_3,ip_12_2,p214,p215);
HA ha46(ip_13_1,ip_14_0,p216,p217);
FA fa62(p164,p166,p168,p218,p219);
HA ha47(p170,p174,p220,p221);
FA fa63(p205,p207,p211,p222,p223);
HA ha48(p213,p215,p224,p225);
FA fa64(p217,p209,p221,p226,p227);
FA fa65(p225,p172,p180,p228,p229);
HA ha49(p219,p223,p230,p231);
FA fa66(p176,p178,p182,p232,p233);
HA ha50(p184,p188,p234,p235);
HA ha51(p227,p231,p236,p237);
HA ha52(p190,p229,p238,p239);
HA ha53(p235,p237,p240,p241);
HA ha54(p186,p233,p242,p243);
HA ha55(p239,p241,p244,p245);
HA ha56(p194,p243,p246,p247);
FA fa67(p245,p192,p247,p248,p249);
FA fa68(p196,p198,p249,p250,p251);
HA ha57(p251,p200,p252,p253);
HA ha58(ip_0_15,ip_1_14,p254,p255);
HA ha59(ip_2_13,ip_3_12,p256,p257);
FA fa69(ip_4_11,ip_5_10,ip_6_9,p258,p259);
HA ha60(ip_7_8,ip_8_7,p260,p261);
HA ha61(ip_9_6,ip_10_5,p262,p263);
FA fa70(ip_11_4,ip_12_3,ip_13_2,p264,p265);
FA fa71(ip_14_1,ip_15_0,p204,p266,p267);
FA fa72(p206,p210,p212,p268,p269);
HA ha62(p214,p216,p270,p271);
HA ha63(p255,p257,p272,p273);
FA fa73(p261,p263,p220,p274,p275);
FA fa74(p224,p259,p265,p276,p277);
HA ha64(p267,p271,p278,p279);
FA fa75(p273,p208,p269,p280,p281);
FA fa76(p275,p279,p218,p282,p283);
HA ha65(p222,p230,p284,p285);
HA ha66(p277,p226,p286,p287);
FA fa77(p234,p236,p281,p288,p289);
FA fa78(p283,p285,p228,p290,p291);
FA fa79(p238,p240,p287,p292,p293);
FA fa80(p232,p242,p244,p294,p295);
HA ha67(p289,p291,p296,p297);
HA ha68(p246,p293,p298,p299);
FA fa81(p297,p295,p299,p300,p301);
FA fa82(p248,p301,p250,p302,p303);
FA fa83(ip_1_15,ip_2_14,ip_3_13,p304,p305);
FA fa84(ip_4_12,ip_5_11,ip_6_10,p306,p307);
FA fa85(ip_7_9,ip_8_8,ip_9_7,p308,p309);
FA fa86(ip_10_6,ip_11_5,ip_12_4,p310,p311);
FA fa87(ip_13_3,ip_14_2,ip_15_1,p312,p313);
FA fa88(p254,p256,p260,p314,p315);
FA fa89(p262,p270,p272,p316,p317);
FA fa90(p305,p307,p309,p318,p319);
FA fa91(p311,p313,p258,p320,p321);
HA ha69(p264,p266,p322,p323);
FA fa92(p278,p315,p268,p324,p325);
FA fa93(p274,p317,p319,p326,p327);
HA ha70(p321,p323,p328,p329);
HA ha71(p276,p284,p330,p331);
HA ha72(p325,p329,p332,p333);
FA fa94(p280,p282,p286,p334,p335);
FA fa95(p327,p331,p333,p336,p337);
FA fa96(p288,p290,p296,p338,p339);
HA ha73(p335,p337,p340,p341);
HA ha74(p292,p298,p342,p343);
FA fa97(p341,p294,p339,p344,p345);
HA ha75(p343,p300,p346,p347);
FA fa98(p345,p347,p302,p348,p349);
FA fa99(ip_2_15,ip_3_14,ip_4_13,p350,p351);
FA fa100(ip_5_12,ip_6_11,ip_7_10,p352,p353);
HA ha76(ip_8_9,ip_9_8,p354,p355);
FA fa101(ip_10_7,ip_11_6,ip_12_5,p356,p357);
HA ha77(ip_13_4,ip_14_3,p358,p359);
FA fa102(ip_15_2,p355,p359,p360,p361);
HA ha78(p351,p353,p362,p363);
HA ha79(p357,p304,p364,p365);
FA fa103(p306,p308,p310,p366,p367);
HA ha80(p312,p361,p368,p369);
HA ha81(p363,p314,p370,p371);
FA fa104(p322,p365,p369,p372,p373);
HA ha82(p316,p318,p374,p375);
FA fa105(p320,p328,p367,p376,p377);
FA fa106(p371,p324,p330,p378,p379);
FA fa107(p332,p373,p375,p380,p381);
HA ha83(p326,p377,p382,p383);
HA ha84(p379,p381,p384,p385);
FA fa108(p383,p334,p336,p386,p387);
HA ha85(p340,p385,p388,p389);
FA fa109(p342,p389,p338,p390,p391);
FA fa110(p387,p391,p344,p392,p393);
HA ha86(p346,p393,p394,p395);
FA fa111(ip_3_15,ip_4_14,ip_5_13,p396,p397);
HA ha87(ip_6_12,ip_7_11,p398,p399);
FA fa112(ip_8_10,ip_9_9,ip_10_8,p400,p401);
HA ha88(ip_11_7,ip_12_6,p402,p403);
HA ha89(ip_13_5,ip_14_4,p404,p405);
HA ha90(ip_15_3,p354,p406,p407);
HA ha91(p358,p399,p408,p409);
FA fa113(p403,p405,p397,p410,p411);
HA ha92(p401,p407,p412,p413);
HA ha93(p409,p350,p414,p415);
FA fa114(p352,p356,p362,p416,p417);
HA ha94(p411,p413,p418,p419);
HA ha95(p360,p364,p420,p421);
HA ha96(p368,p415,p422,p423);
FA fa115(p419,p370,p417,p424,p425);
HA ha97(p421,p423,p426,p427);
FA fa116(p366,p374,p427,p428,p429);
HA ha98(p372,p425,p430,p431);
HA ha99(p376,p382,p432,p433);
FA fa117(p429,p431,p378,p434,p435);
FA fa118(p380,p384,p433,p436,p437);
HA ha100(p388,p435,p438,p439);
FA fa119(p437,p439,p386,p440,p441);
FA fa120(p390,p441,p392,p442,p443);
HA ha101(ip_4_15,ip_5_14,p444,p445);
HA ha102(ip_6_13,ip_7_12,p446,p447);
FA fa121(ip_8_11,ip_9_10,ip_10_9,p448,p449);
HA ha103(ip_11_8,ip_12_7,p450,p451);
FA fa122(ip_13_6,ip_14_5,ip_15_4,p452,p453);
HA ha104(p398,p402,p454,p455);
HA ha105(p404,p445,p456,p457);
FA fa123(p447,p451,p406,p458,p459);
FA fa124(p408,p449,p453,p460,p461);
HA ha106(p455,p457,p462,p463);
HA ha107(p396,p400,p464,p465);
HA ha108(p412,p459,p466,p467);
HA ha109(p463,p410,p468,p469);
FA fa125(p414,p418,p461,p470,p471);
HA ha110(p465,p467,p472,p473);
HA ha111(p420,p422,p474,p475);
HA ha112(p469,p473,p476,p477);
FA fa126(p416,p426,p471,p478,p479);
HA ha113(p475,p477,p480,p481);
FA fa127(p481,p424,p430,p482,p483);
FA fa128(p479,p428,p432,p484,p485);
FA fa129(p483,p434,p438,p486,p487);
FA fa130(p485,p436,p487,p488,p489);
HA ha114(p440,p489,p490,p491);
FA fa131(ip_5_15,ip_6_14,ip_7_13,p492,p493);
FA fa132(ip_8_12,ip_9_11,ip_10_10,p494,p495);
FA fa133(ip_11_9,ip_12_8,ip_13_7,p496,p497);
FA fa134(ip_14_6,ip_15_5,p444,p498,p499);
FA fa135(p446,p450,p454,p500,p501);
FA fa136(p456,p493,p495,p502,p503);
HA ha115(p497,p499,p504,p505);
FA fa137(p448,p452,p462,p506,p507);
HA ha116(p501,p505,p508,p509);
FA fa138(p458,p464,p466,p510,p511);
HA ha117(p503,p509,p512,p513);
HA ha118(p460,p468,p514,p515);
HA ha119(p472,p507,p516,p517);
FA fa139(p513,p474,p476,p518,p519);
HA ha120(p511,p515,p520,p521);
HA ha121(p517,p470,p522,p523);
FA fa140(p480,p521,p519,p524,p525);
HA ha122(p523,p478,p526,p527);
HA ha123(p525,p527,p528,p529);
FA fa141(p482,p529,p484,p530,p531);
FA fa142(p531,p486,p488,p532,p533);
FA fa143(ip_6_15,ip_7_14,ip_8_13,p534,p535);
HA ha124(ip_9_12,ip_10_11,p536,p537);
FA fa144(ip_11_10,ip_12_9,ip_13_8,p538,p539);
HA ha125(ip_14_7,ip_15_6,p540,p541);
FA fa145(p537,p541,p535,p542,p543);
FA fa146(p539,p492,p494,p544,p545);
FA fa147(p496,p498,p504,p546,p547);
HA ha126(p543,p500,p548,p549);
FA fa148(p508,p502,p512,p550,p551);
HA ha127(p545,p547,p552,p553);
FA fa149(p549,p506,p514,p554,p555);
FA fa150(p516,p553,p510,p556,p557);
HA ha128(p520,p551,p558,p559);
HA ha129(p522,p555,p560,p561);
HA ha130(p557,p559,p562,p563);
HA ha131(p518,p561,p564,p565);
FA fa151(p563,p524,p526,p566,p567);
FA fa152(p565,p528,p567,p568,p569);
FA fa153(p569,p530,p532,p570,p571);
HA ha132(ip_7_15,ip_8_14,p572,p573);
HA ha133(ip_9_13,ip_10_12,p574,p575);
HA ha134(ip_11_11,ip_12_10,p576,p577);
HA ha135(ip_13_9,ip_14_8,p578,p579);
FA fa154(ip_15_7,p536,p540,p580,p581);
FA fa155(p573,p575,p577,p582,p583);
HA ha136(p579,p534,p584,p585);
HA ha137(p538,p581,p586,p587);
HA ha138(p583,p542,p588,p589);
FA fa156(p585,p587,p548,p590,p591);
FA fa157(p589,p544,p546,p592,p593);
HA ha139(p552,p591,p594,p595);
HA ha140(p595,p550,p596,p597);
FA fa158(p558,p593,p554,p598,p599);
FA fa159(p556,p560,p562,p600,p601);
HA ha141(p597,p564,p602,p603);
HA ha142(p599,p601,p604,p605);
FA fa160(p603,p605,p566,p606,p607);
FA fa161(p568,p607,p570,p608,p609);
HA ha143(ip_8_15,ip_9_14,p610,p611);
FA fa162(ip_10_13,ip_11_12,ip_12_11,p612,p613);
HA ha144(ip_13_10,ip_14_9,p614,p615);
FA fa163(ip_15_8,p572,p574,p616,p617);
FA fa164(p576,p578,p611,p618,p619);
HA ha145(p615,p613,p620,p621);
FA fa165(p617,p619,p621,p622,p623);
FA fa166(p580,p582,p584,p624,p625);
HA ha146(p586,p588,p626,p627);
FA fa167(p623,p625,p627,p628,p629);
FA fa168(p590,p594,p629,p630,p631);
FA fa169(p592,p596,p631,p632,p633);
HA ha147(p598,p602,p634,p635);
HA ha148(p633,p600,p636,p637);
FA fa170(p604,p635,p637,p638,p639);
HA ha149(p639,p606,p640,p641);
FA fa171(ip_9_15,ip_10_14,ip_11_13,p642,p643);
FA fa172(ip_12_12,ip_13_11,ip_14_10,p644,p645);
FA fa173(ip_15_9,p610,p614,p646,p647);
HA ha150(p643,p645,p648,p649);
FA fa174(p612,p620,p647,p650,p651);
FA fa175(p649,p616,p618,p652,p653);
FA fa176(p651,p622,p626,p654,p655);
FA fa177(p653,p624,p655,p656,p657);
HA ha151(p628,p657,p658,p659);
HA ha152(p630,p659,p660,p661);
FA fa178(p661,p632,p634,p662,p663);
HA ha153(p636,p663,p664,p665);
HA ha154(p638,p665,p666,p667);
FA fa179(ip_10_15,ip_11_14,ip_12_13,p668,p669);
FA fa180(ip_13_12,ip_14_11,ip_15_10,p670,p671);
HA ha155(p669,p671,p672,p673);
HA ha156(p642,p644,p674,p675);
HA ha157(p648,p673,p676,p677);
HA ha158(p646,p675,p678,p679);
FA fa181(p677,p679,p650,p680,p681);
FA fa182(p652,p681,p654,p682,p683);
HA ha159(p656,p658,p684,p685);
HA ha160(p683,p660,p686,p687);
HA ha161(p685,p687,p688,p689);
HA ha162(p689,p662,p690,p691);
HA ha163(p664,p666,p692,p693);
FA fa183(ip_11_15,ip_12_14,ip_13_13,p694,p695);
FA fa184(ip_14_12,ip_15_11,p695,p696,p697);
FA fa185(p668,p670,p672,p698,p699);
HA ha164(p697,p674,p700,p701);
HA ha165(p676,p678,p702,p703);
HA ha166(p699,p701,p704,p705);
FA fa186(p703,p705,p680,p706,p707);
FA fa187(p707,p682,p684,p708,p709);
FA fa188(p686,p688,p709,p710,p711);
FA fa189(p711,p690,p692,p712,p713);
FA fa190(ip_12_15,ip_13_14,ip_14_13,p714,p715);
HA ha167(ip_15_12,p715,p716,p717);
FA fa191(p694,p717,p696,p718,p719);
HA ha168(p700,p719,p720,p721);
HA ha169(p698,p702,p722,p723);
FA fa192(p704,p721,p723,p724,p725);
FA fa193(p725,p706,p708,p726,p727);
FA fa194(p727,p710,p712,p728,p729);
FA fa195(ip_13_15,ip_14_14,ip_15_13,p730,p731);
FA fa196(p731,p714,p716,p732,p733);
FA fa197(p733,p718,p720,p734,p735);
HA ha170(p722,p735,p736,p737);
HA ha171(p724,p737,p738,p739);
FA fa198(p739,p726,p728,p740,p741);
FA fa199(ip_14_15,ip_15_14,p730,p742,p743);
FA fa200(p743,p732,p734,p744,p745);
FA fa201(p736,p738,p745,p746,p747);
FA fa202(ip_15_15,p742,p744,p748,p749);
wire [31:0] a,b;
wire [31:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p5;
assign b[3] = 1'b0;
assign a[4] = p11;
assign b[4] = p4;
assign a[5] = p10;
assign b[5] = p19;
assign a[6] = p18;
assign b[6] = p29;
assign a[7] = p28;
assign b[7] = p43;
assign a[8] = p59;
assign b[8] = 1'b0;
assign a[9] = p79;
assign b[9] = p58;
assign a[10] = p78;
assign b[10] = p103;
assign a[11] = p102;
assign b[11] = p133;
assign a[12] = p161;
assign b[12] = p163;
assign a[13] = p162;
assign b[13] = p203;
assign a[14] = p202;
assign b[14] = p253;
assign a[15] = p252;
assign b[15] = p303;
assign a[16] = p349;
assign b[16] = 1'b0;
assign a[17] = p395;
assign b[17] = p348;
assign a[18] = p394;
assign b[18] = p443;
assign a[19] = p491;
assign b[19] = p442;
assign a[20] = p490;
assign b[20] = p533;
assign a[21] = p571;
assign b[21] = 1'b0;
assign a[22] = p609;
assign b[22] = 1'b0;
assign a[23] = p641;
assign b[23] = p608;
assign a[24] = p640;
assign b[24] = p667;
assign a[25] = p691;
assign b[25] = p693;
assign a[26] = p713;
assign b[26] = 1'b0;
assign a[27] = p729;
assign b[27] = 1'b0;
assign a[28] = p741;
assign b[28] = 1'b0;
assign a[29] = p747;
assign b[29] = p740;
assign a[30] = p749;
assign b[30] = p746;
assign a[31] = p748;
assign b[31] = 1'b0;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[31] = s[31];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [31:0] a,b;
output [31:0] s;
assign s = a+b;
endmodule
