// 1 2 2 2 2 2 2 2 1 2 1 1 1 2 1 2 2 2 1 2 2 1 2 1 2 2 2 1 2 1 1 1 2 2 2 2 2 1 2 1 2 2 1 2 2 1 2 2 1 1 1 1 2 2 2 1 1 1 2 1 2 1 1 1 1 1 2 2 2 1 1 1 1 2 2 1 2 1 2 1 2 2 2 2 2 2 2 2 1 1 2 2 1 1 2 1 2 1 2 2 2 1 2 2 2 2 1 2 2 1 2 1 2 1 2 2 1 1 1 1 1 2 1 1 2 1 2 1 

module main(x,y,o);
input [63:0] x,y;
output [127:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_0_16,ip_0_17,ip_0_18,ip_0_19,ip_0_20,ip_0_21,ip_0_22,ip_0_23,ip_0_24,ip_0_25,ip_0_26,ip_0_27,ip_0_28,ip_0_29,ip_0_30,ip_0_31,ip_0_32,ip_0_33,ip_0_34,ip_0_35,ip_0_36,ip_0_37,ip_0_38,ip_0_39,ip_0_40,ip_0_41,ip_0_42,ip_0_43,ip_0_44,ip_0_45,ip_0_46,ip_0_47,ip_0_48,ip_0_49,ip_0_50,ip_0_51,ip_0_52,ip_0_53,ip_0_54,ip_0_55,ip_0_56,ip_0_57,ip_0_58,ip_0_59,ip_0_60,ip_0_61,ip_0_62,ip_0_63,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_1_16,ip_1_17,ip_1_18,ip_1_19,ip_1_20,ip_1_21,ip_1_22,ip_1_23,ip_1_24,ip_1_25,ip_1_26,ip_1_27,ip_1_28,ip_1_29,ip_1_30,ip_1_31,ip_1_32,ip_1_33,ip_1_34,ip_1_35,ip_1_36,ip_1_37,ip_1_38,ip_1_39,ip_1_40,ip_1_41,ip_1_42,ip_1_43,ip_1_44,ip_1_45,ip_1_46,ip_1_47,ip_1_48,ip_1_49,ip_1_50,ip_1_51,ip_1_52,ip_1_53,ip_1_54,ip_1_55,ip_1_56,ip_1_57,ip_1_58,ip_1_59,ip_1_60,ip_1_61,ip_1_62,ip_1_63,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_2_16,ip_2_17,ip_2_18,ip_2_19,ip_2_20,ip_2_21,ip_2_22,ip_2_23,ip_2_24,ip_2_25,ip_2_26,ip_2_27,ip_2_28,ip_2_29,ip_2_30,ip_2_31,ip_2_32,ip_2_33,ip_2_34,ip_2_35,ip_2_36,ip_2_37,ip_2_38,ip_2_39,ip_2_40,ip_2_41,ip_2_42,ip_2_43,ip_2_44,ip_2_45,ip_2_46,ip_2_47,ip_2_48,ip_2_49,ip_2_50,ip_2_51,ip_2_52,ip_2_53,ip_2_54,ip_2_55,ip_2_56,ip_2_57,ip_2_58,ip_2_59,ip_2_60,ip_2_61,ip_2_62,ip_2_63,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_3_16,ip_3_17,ip_3_18,ip_3_19,ip_3_20,ip_3_21,ip_3_22,ip_3_23,ip_3_24,ip_3_25,ip_3_26,ip_3_27,ip_3_28,ip_3_29,ip_3_30,ip_3_31,ip_3_32,ip_3_33,ip_3_34,ip_3_35,ip_3_36,ip_3_37,ip_3_38,ip_3_39,ip_3_40,ip_3_41,ip_3_42,ip_3_43,ip_3_44,ip_3_45,ip_3_46,ip_3_47,ip_3_48,ip_3_49,ip_3_50,ip_3_51,ip_3_52,ip_3_53,ip_3_54,ip_3_55,ip_3_56,ip_3_57,ip_3_58,ip_3_59,ip_3_60,ip_3_61,ip_3_62,ip_3_63,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_4_16,ip_4_17,ip_4_18,ip_4_19,ip_4_20,ip_4_21,ip_4_22,ip_4_23,ip_4_24,ip_4_25,ip_4_26,ip_4_27,ip_4_28,ip_4_29,ip_4_30,ip_4_31,ip_4_32,ip_4_33,ip_4_34,ip_4_35,ip_4_36,ip_4_37,ip_4_38,ip_4_39,ip_4_40,ip_4_41,ip_4_42,ip_4_43,ip_4_44,ip_4_45,ip_4_46,ip_4_47,ip_4_48,ip_4_49,ip_4_50,ip_4_51,ip_4_52,ip_4_53,ip_4_54,ip_4_55,ip_4_56,ip_4_57,ip_4_58,ip_4_59,ip_4_60,ip_4_61,ip_4_62,ip_4_63,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_5_16,ip_5_17,ip_5_18,ip_5_19,ip_5_20,ip_5_21,ip_5_22,ip_5_23,ip_5_24,ip_5_25,ip_5_26,ip_5_27,ip_5_28,ip_5_29,ip_5_30,ip_5_31,ip_5_32,ip_5_33,ip_5_34,ip_5_35,ip_5_36,ip_5_37,ip_5_38,ip_5_39,ip_5_40,ip_5_41,ip_5_42,ip_5_43,ip_5_44,ip_5_45,ip_5_46,ip_5_47,ip_5_48,ip_5_49,ip_5_50,ip_5_51,ip_5_52,ip_5_53,ip_5_54,ip_5_55,ip_5_56,ip_5_57,ip_5_58,ip_5_59,ip_5_60,ip_5_61,ip_5_62,ip_5_63,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_6_16,ip_6_17,ip_6_18,ip_6_19,ip_6_20,ip_6_21,ip_6_22,ip_6_23,ip_6_24,ip_6_25,ip_6_26,ip_6_27,ip_6_28,ip_6_29,ip_6_30,ip_6_31,ip_6_32,ip_6_33,ip_6_34,ip_6_35,ip_6_36,ip_6_37,ip_6_38,ip_6_39,ip_6_40,ip_6_41,ip_6_42,ip_6_43,ip_6_44,ip_6_45,ip_6_46,ip_6_47,ip_6_48,ip_6_49,ip_6_50,ip_6_51,ip_6_52,ip_6_53,ip_6_54,ip_6_55,ip_6_56,ip_6_57,ip_6_58,ip_6_59,ip_6_60,ip_6_61,ip_6_62,ip_6_63,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_7_16,ip_7_17,ip_7_18,ip_7_19,ip_7_20,ip_7_21,ip_7_22,ip_7_23,ip_7_24,ip_7_25,ip_7_26,ip_7_27,ip_7_28,ip_7_29,ip_7_30,ip_7_31,ip_7_32,ip_7_33,ip_7_34,ip_7_35,ip_7_36,ip_7_37,ip_7_38,ip_7_39,ip_7_40,ip_7_41,ip_7_42,ip_7_43,ip_7_44,ip_7_45,ip_7_46,ip_7_47,ip_7_48,ip_7_49,ip_7_50,ip_7_51,ip_7_52,ip_7_53,ip_7_54,ip_7_55,ip_7_56,ip_7_57,ip_7_58,ip_7_59,ip_7_60,ip_7_61,ip_7_62,ip_7_63,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_8_16,ip_8_17,ip_8_18,ip_8_19,ip_8_20,ip_8_21,ip_8_22,ip_8_23,ip_8_24,ip_8_25,ip_8_26,ip_8_27,ip_8_28,ip_8_29,ip_8_30,ip_8_31,ip_8_32,ip_8_33,ip_8_34,ip_8_35,ip_8_36,ip_8_37,ip_8_38,ip_8_39,ip_8_40,ip_8_41,ip_8_42,ip_8_43,ip_8_44,ip_8_45,ip_8_46,ip_8_47,ip_8_48,ip_8_49,ip_8_50,ip_8_51,ip_8_52,ip_8_53,ip_8_54,ip_8_55,ip_8_56,ip_8_57,ip_8_58,ip_8_59,ip_8_60,ip_8_61,ip_8_62,ip_8_63,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_9_16,ip_9_17,ip_9_18,ip_9_19,ip_9_20,ip_9_21,ip_9_22,ip_9_23,ip_9_24,ip_9_25,ip_9_26,ip_9_27,ip_9_28,ip_9_29,ip_9_30,ip_9_31,ip_9_32,ip_9_33,ip_9_34,ip_9_35,ip_9_36,ip_9_37,ip_9_38,ip_9_39,ip_9_40,ip_9_41,ip_9_42,ip_9_43,ip_9_44,ip_9_45,ip_9_46,ip_9_47,ip_9_48,ip_9_49,ip_9_50,ip_9_51,ip_9_52,ip_9_53,ip_9_54,ip_9_55,ip_9_56,ip_9_57,ip_9_58,ip_9_59,ip_9_60,ip_9_61,ip_9_62,ip_9_63,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_10_16,ip_10_17,ip_10_18,ip_10_19,ip_10_20,ip_10_21,ip_10_22,ip_10_23,ip_10_24,ip_10_25,ip_10_26,ip_10_27,ip_10_28,ip_10_29,ip_10_30,ip_10_31,ip_10_32,ip_10_33,ip_10_34,ip_10_35,ip_10_36,ip_10_37,ip_10_38,ip_10_39,ip_10_40,ip_10_41,ip_10_42,ip_10_43,ip_10_44,ip_10_45,ip_10_46,ip_10_47,ip_10_48,ip_10_49,ip_10_50,ip_10_51,ip_10_52,ip_10_53,ip_10_54,ip_10_55,ip_10_56,ip_10_57,ip_10_58,ip_10_59,ip_10_60,ip_10_61,ip_10_62,ip_10_63,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_11_16,ip_11_17,ip_11_18,ip_11_19,ip_11_20,ip_11_21,ip_11_22,ip_11_23,ip_11_24,ip_11_25,ip_11_26,ip_11_27,ip_11_28,ip_11_29,ip_11_30,ip_11_31,ip_11_32,ip_11_33,ip_11_34,ip_11_35,ip_11_36,ip_11_37,ip_11_38,ip_11_39,ip_11_40,ip_11_41,ip_11_42,ip_11_43,ip_11_44,ip_11_45,ip_11_46,ip_11_47,ip_11_48,ip_11_49,ip_11_50,ip_11_51,ip_11_52,ip_11_53,ip_11_54,ip_11_55,ip_11_56,ip_11_57,ip_11_58,ip_11_59,ip_11_60,ip_11_61,ip_11_62,ip_11_63,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_12_16,ip_12_17,ip_12_18,ip_12_19,ip_12_20,ip_12_21,ip_12_22,ip_12_23,ip_12_24,ip_12_25,ip_12_26,ip_12_27,ip_12_28,ip_12_29,ip_12_30,ip_12_31,ip_12_32,ip_12_33,ip_12_34,ip_12_35,ip_12_36,ip_12_37,ip_12_38,ip_12_39,ip_12_40,ip_12_41,ip_12_42,ip_12_43,ip_12_44,ip_12_45,ip_12_46,ip_12_47,ip_12_48,ip_12_49,ip_12_50,ip_12_51,ip_12_52,ip_12_53,ip_12_54,ip_12_55,ip_12_56,ip_12_57,ip_12_58,ip_12_59,ip_12_60,ip_12_61,ip_12_62,ip_12_63,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_13_16,ip_13_17,ip_13_18,ip_13_19,ip_13_20,ip_13_21,ip_13_22,ip_13_23,ip_13_24,ip_13_25,ip_13_26,ip_13_27,ip_13_28,ip_13_29,ip_13_30,ip_13_31,ip_13_32,ip_13_33,ip_13_34,ip_13_35,ip_13_36,ip_13_37,ip_13_38,ip_13_39,ip_13_40,ip_13_41,ip_13_42,ip_13_43,ip_13_44,ip_13_45,ip_13_46,ip_13_47,ip_13_48,ip_13_49,ip_13_50,ip_13_51,ip_13_52,ip_13_53,ip_13_54,ip_13_55,ip_13_56,ip_13_57,ip_13_58,ip_13_59,ip_13_60,ip_13_61,ip_13_62,ip_13_63,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_14_16,ip_14_17,ip_14_18,ip_14_19,ip_14_20,ip_14_21,ip_14_22,ip_14_23,ip_14_24,ip_14_25,ip_14_26,ip_14_27,ip_14_28,ip_14_29,ip_14_30,ip_14_31,ip_14_32,ip_14_33,ip_14_34,ip_14_35,ip_14_36,ip_14_37,ip_14_38,ip_14_39,ip_14_40,ip_14_41,ip_14_42,ip_14_43,ip_14_44,ip_14_45,ip_14_46,ip_14_47,ip_14_48,ip_14_49,ip_14_50,ip_14_51,ip_14_52,ip_14_53,ip_14_54,ip_14_55,ip_14_56,ip_14_57,ip_14_58,ip_14_59,ip_14_60,ip_14_61,ip_14_62,ip_14_63,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15,ip_15_16,ip_15_17,ip_15_18,ip_15_19,ip_15_20,ip_15_21,ip_15_22,ip_15_23,ip_15_24,ip_15_25,ip_15_26,ip_15_27,ip_15_28,ip_15_29,ip_15_30,ip_15_31,ip_15_32,ip_15_33,ip_15_34,ip_15_35,ip_15_36,ip_15_37,ip_15_38,ip_15_39,ip_15_40,ip_15_41,ip_15_42,ip_15_43,ip_15_44,ip_15_45,ip_15_46,ip_15_47,ip_15_48,ip_15_49,ip_15_50,ip_15_51,ip_15_52,ip_15_53,ip_15_54,ip_15_55,ip_15_56,ip_15_57,ip_15_58,ip_15_59,ip_15_60,ip_15_61,ip_15_62,ip_15_63,ip_16_0,ip_16_1,ip_16_2,ip_16_3,ip_16_4,ip_16_5,ip_16_6,ip_16_7,ip_16_8,ip_16_9,ip_16_10,ip_16_11,ip_16_12,ip_16_13,ip_16_14,ip_16_15,ip_16_16,ip_16_17,ip_16_18,ip_16_19,ip_16_20,ip_16_21,ip_16_22,ip_16_23,ip_16_24,ip_16_25,ip_16_26,ip_16_27,ip_16_28,ip_16_29,ip_16_30,ip_16_31,ip_16_32,ip_16_33,ip_16_34,ip_16_35,ip_16_36,ip_16_37,ip_16_38,ip_16_39,ip_16_40,ip_16_41,ip_16_42,ip_16_43,ip_16_44,ip_16_45,ip_16_46,ip_16_47,ip_16_48,ip_16_49,ip_16_50,ip_16_51,ip_16_52,ip_16_53,ip_16_54,ip_16_55,ip_16_56,ip_16_57,ip_16_58,ip_16_59,ip_16_60,ip_16_61,ip_16_62,ip_16_63,ip_17_0,ip_17_1,ip_17_2,ip_17_3,ip_17_4,ip_17_5,ip_17_6,ip_17_7,ip_17_8,ip_17_9,ip_17_10,ip_17_11,ip_17_12,ip_17_13,ip_17_14,ip_17_15,ip_17_16,ip_17_17,ip_17_18,ip_17_19,ip_17_20,ip_17_21,ip_17_22,ip_17_23,ip_17_24,ip_17_25,ip_17_26,ip_17_27,ip_17_28,ip_17_29,ip_17_30,ip_17_31,ip_17_32,ip_17_33,ip_17_34,ip_17_35,ip_17_36,ip_17_37,ip_17_38,ip_17_39,ip_17_40,ip_17_41,ip_17_42,ip_17_43,ip_17_44,ip_17_45,ip_17_46,ip_17_47,ip_17_48,ip_17_49,ip_17_50,ip_17_51,ip_17_52,ip_17_53,ip_17_54,ip_17_55,ip_17_56,ip_17_57,ip_17_58,ip_17_59,ip_17_60,ip_17_61,ip_17_62,ip_17_63,ip_18_0,ip_18_1,ip_18_2,ip_18_3,ip_18_4,ip_18_5,ip_18_6,ip_18_7,ip_18_8,ip_18_9,ip_18_10,ip_18_11,ip_18_12,ip_18_13,ip_18_14,ip_18_15,ip_18_16,ip_18_17,ip_18_18,ip_18_19,ip_18_20,ip_18_21,ip_18_22,ip_18_23,ip_18_24,ip_18_25,ip_18_26,ip_18_27,ip_18_28,ip_18_29,ip_18_30,ip_18_31,ip_18_32,ip_18_33,ip_18_34,ip_18_35,ip_18_36,ip_18_37,ip_18_38,ip_18_39,ip_18_40,ip_18_41,ip_18_42,ip_18_43,ip_18_44,ip_18_45,ip_18_46,ip_18_47,ip_18_48,ip_18_49,ip_18_50,ip_18_51,ip_18_52,ip_18_53,ip_18_54,ip_18_55,ip_18_56,ip_18_57,ip_18_58,ip_18_59,ip_18_60,ip_18_61,ip_18_62,ip_18_63,ip_19_0,ip_19_1,ip_19_2,ip_19_3,ip_19_4,ip_19_5,ip_19_6,ip_19_7,ip_19_8,ip_19_9,ip_19_10,ip_19_11,ip_19_12,ip_19_13,ip_19_14,ip_19_15,ip_19_16,ip_19_17,ip_19_18,ip_19_19,ip_19_20,ip_19_21,ip_19_22,ip_19_23,ip_19_24,ip_19_25,ip_19_26,ip_19_27,ip_19_28,ip_19_29,ip_19_30,ip_19_31,ip_19_32,ip_19_33,ip_19_34,ip_19_35,ip_19_36,ip_19_37,ip_19_38,ip_19_39,ip_19_40,ip_19_41,ip_19_42,ip_19_43,ip_19_44,ip_19_45,ip_19_46,ip_19_47,ip_19_48,ip_19_49,ip_19_50,ip_19_51,ip_19_52,ip_19_53,ip_19_54,ip_19_55,ip_19_56,ip_19_57,ip_19_58,ip_19_59,ip_19_60,ip_19_61,ip_19_62,ip_19_63,ip_20_0,ip_20_1,ip_20_2,ip_20_3,ip_20_4,ip_20_5,ip_20_6,ip_20_7,ip_20_8,ip_20_9,ip_20_10,ip_20_11,ip_20_12,ip_20_13,ip_20_14,ip_20_15,ip_20_16,ip_20_17,ip_20_18,ip_20_19,ip_20_20,ip_20_21,ip_20_22,ip_20_23,ip_20_24,ip_20_25,ip_20_26,ip_20_27,ip_20_28,ip_20_29,ip_20_30,ip_20_31,ip_20_32,ip_20_33,ip_20_34,ip_20_35,ip_20_36,ip_20_37,ip_20_38,ip_20_39,ip_20_40,ip_20_41,ip_20_42,ip_20_43,ip_20_44,ip_20_45,ip_20_46,ip_20_47,ip_20_48,ip_20_49,ip_20_50,ip_20_51,ip_20_52,ip_20_53,ip_20_54,ip_20_55,ip_20_56,ip_20_57,ip_20_58,ip_20_59,ip_20_60,ip_20_61,ip_20_62,ip_20_63,ip_21_0,ip_21_1,ip_21_2,ip_21_3,ip_21_4,ip_21_5,ip_21_6,ip_21_7,ip_21_8,ip_21_9,ip_21_10,ip_21_11,ip_21_12,ip_21_13,ip_21_14,ip_21_15,ip_21_16,ip_21_17,ip_21_18,ip_21_19,ip_21_20,ip_21_21,ip_21_22,ip_21_23,ip_21_24,ip_21_25,ip_21_26,ip_21_27,ip_21_28,ip_21_29,ip_21_30,ip_21_31,ip_21_32,ip_21_33,ip_21_34,ip_21_35,ip_21_36,ip_21_37,ip_21_38,ip_21_39,ip_21_40,ip_21_41,ip_21_42,ip_21_43,ip_21_44,ip_21_45,ip_21_46,ip_21_47,ip_21_48,ip_21_49,ip_21_50,ip_21_51,ip_21_52,ip_21_53,ip_21_54,ip_21_55,ip_21_56,ip_21_57,ip_21_58,ip_21_59,ip_21_60,ip_21_61,ip_21_62,ip_21_63,ip_22_0,ip_22_1,ip_22_2,ip_22_3,ip_22_4,ip_22_5,ip_22_6,ip_22_7,ip_22_8,ip_22_9,ip_22_10,ip_22_11,ip_22_12,ip_22_13,ip_22_14,ip_22_15,ip_22_16,ip_22_17,ip_22_18,ip_22_19,ip_22_20,ip_22_21,ip_22_22,ip_22_23,ip_22_24,ip_22_25,ip_22_26,ip_22_27,ip_22_28,ip_22_29,ip_22_30,ip_22_31,ip_22_32,ip_22_33,ip_22_34,ip_22_35,ip_22_36,ip_22_37,ip_22_38,ip_22_39,ip_22_40,ip_22_41,ip_22_42,ip_22_43,ip_22_44,ip_22_45,ip_22_46,ip_22_47,ip_22_48,ip_22_49,ip_22_50,ip_22_51,ip_22_52,ip_22_53,ip_22_54,ip_22_55,ip_22_56,ip_22_57,ip_22_58,ip_22_59,ip_22_60,ip_22_61,ip_22_62,ip_22_63,ip_23_0,ip_23_1,ip_23_2,ip_23_3,ip_23_4,ip_23_5,ip_23_6,ip_23_7,ip_23_8,ip_23_9,ip_23_10,ip_23_11,ip_23_12,ip_23_13,ip_23_14,ip_23_15,ip_23_16,ip_23_17,ip_23_18,ip_23_19,ip_23_20,ip_23_21,ip_23_22,ip_23_23,ip_23_24,ip_23_25,ip_23_26,ip_23_27,ip_23_28,ip_23_29,ip_23_30,ip_23_31,ip_23_32,ip_23_33,ip_23_34,ip_23_35,ip_23_36,ip_23_37,ip_23_38,ip_23_39,ip_23_40,ip_23_41,ip_23_42,ip_23_43,ip_23_44,ip_23_45,ip_23_46,ip_23_47,ip_23_48,ip_23_49,ip_23_50,ip_23_51,ip_23_52,ip_23_53,ip_23_54,ip_23_55,ip_23_56,ip_23_57,ip_23_58,ip_23_59,ip_23_60,ip_23_61,ip_23_62,ip_23_63,ip_24_0,ip_24_1,ip_24_2,ip_24_3,ip_24_4,ip_24_5,ip_24_6,ip_24_7,ip_24_8,ip_24_9,ip_24_10,ip_24_11,ip_24_12,ip_24_13,ip_24_14,ip_24_15,ip_24_16,ip_24_17,ip_24_18,ip_24_19,ip_24_20,ip_24_21,ip_24_22,ip_24_23,ip_24_24,ip_24_25,ip_24_26,ip_24_27,ip_24_28,ip_24_29,ip_24_30,ip_24_31,ip_24_32,ip_24_33,ip_24_34,ip_24_35,ip_24_36,ip_24_37,ip_24_38,ip_24_39,ip_24_40,ip_24_41,ip_24_42,ip_24_43,ip_24_44,ip_24_45,ip_24_46,ip_24_47,ip_24_48,ip_24_49,ip_24_50,ip_24_51,ip_24_52,ip_24_53,ip_24_54,ip_24_55,ip_24_56,ip_24_57,ip_24_58,ip_24_59,ip_24_60,ip_24_61,ip_24_62,ip_24_63,ip_25_0,ip_25_1,ip_25_2,ip_25_3,ip_25_4,ip_25_5,ip_25_6,ip_25_7,ip_25_8,ip_25_9,ip_25_10,ip_25_11,ip_25_12,ip_25_13,ip_25_14,ip_25_15,ip_25_16,ip_25_17,ip_25_18,ip_25_19,ip_25_20,ip_25_21,ip_25_22,ip_25_23,ip_25_24,ip_25_25,ip_25_26,ip_25_27,ip_25_28,ip_25_29,ip_25_30,ip_25_31,ip_25_32,ip_25_33,ip_25_34,ip_25_35,ip_25_36,ip_25_37,ip_25_38,ip_25_39,ip_25_40,ip_25_41,ip_25_42,ip_25_43,ip_25_44,ip_25_45,ip_25_46,ip_25_47,ip_25_48,ip_25_49,ip_25_50,ip_25_51,ip_25_52,ip_25_53,ip_25_54,ip_25_55,ip_25_56,ip_25_57,ip_25_58,ip_25_59,ip_25_60,ip_25_61,ip_25_62,ip_25_63,ip_26_0,ip_26_1,ip_26_2,ip_26_3,ip_26_4,ip_26_5,ip_26_6,ip_26_7,ip_26_8,ip_26_9,ip_26_10,ip_26_11,ip_26_12,ip_26_13,ip_26_14,ip_26_15,ip_26_16,ip_26_17,ip_26_18,ip_26_19,ip_26_20,ip_26_21,ip_26_22,ip_26_23,ip_26_24,ip_26_25,ip_26_26,ip_26_27,ip_26_28,ip_26_29,ip_26_30,ip_26_31,ip_26_32,ip_26_33,ip_26_34,ip_26_35,ip_26_36,ip_26_37,ip_26_38,ip_26_39,ip_26_40,ip_26_41,ip_26_42,ip_26_43,ip_26_44,ip_26_45,ip_26_46,ip_26_47,ip_26_48,ip_26_49,ip_26_50,ip_26_51,ip_26_52,ip_26_53,ip_26_54,ip_26_55,ip_26_56,ip_26_57,ip_26_58,ip_26_59,ip_26_60,ip_26_61,ip_26_62,ip_26_63,ip_27_0,ip_27_1,ip_27_2,ip_27_3,ip_27_4,ip_27_5,ip_27_6,ip_27_7,ip_27_8,ip_27_9,ip_27_10,ip_27_11,ip_27_12,ip_27_13,ip_27_14,ip_27_15,ip_27_16,ip_27_17,ip_27_18,ip_27_19,ip_27_20,ip_27_21,ip_27_22,ip_27_23,ip_27_24,ip_27_25,ip_27_26,ip_27_27,ip_27_28,ip_27_29,ip_27_30,ip_27_31,ip_27_32,ip_27_33,ip_27_34,ip_27_35,ip_27_36,ip_27_37,ip_27_38,ip_27_39,ip_27_40,ip_27_41,ip_27_42,ip_27_43,ip_27_44,ip_27_45,ip_27_46,ip_27_47,ip_27_48,ip_27_49,ip_27_50,ip_27_51,ip_27_52,ip_27_53,ip_27_54,ip_27_55,ip_27_56,ip_27_57,ip_27_58,ip_27_59,ip_27_60,ip_27_61,ip_27_62,ip_27_63,ip_28_0,ip_28_1,ip_28_2,ip_28_3,ip_28_4,ip_28_5,ip_28_6,ip_28_7,ip_28_8,ip_28_9,ip_28_10,ip_28_11,ip_28_12,ip_28_13,ip_28_14,ip_28_15,ip_28_16,ip_28_17,ip_28_18,ip_28_19,ip_28_20,ip_28_21,ip_28_22,ip_28_23,ip_28_24,ip_28_25,ip_28_26,ip_28_27,ip_28_28,ip_28_29,ip_28_30,ip_28_31,ip_28_32,ip_28_33,ip_28_34,ip_28_35,ip_28_36,ip_28_37,ip_28_38,ip_28_39,ip_28_40,ip_28_41,ip_28_42,ip_28_43,ip_28_44,ip_28_45,ip_28_46,ip_28_47,ip_28_48,ip_28_49,ip_28_50,ip_28_51,ip_28_52,ip_28_53,ip_28_54,ip_28_55,ip_28_56,ip_28_57,ip_28_58,ip_28_59,ip_28_60,ip_28_61,ip_28_62,ip_28_63,ip_29_0,ip_29_1,ip_29_2,ip_29_3,ip_29_4,ip_29_5,ip_29_6,ip_29_7,ip_29_8,ip_29_9,ip_29_10,ip_29_11,ip_29_12,ip_29_13,ip_29_14,ip_29_15,ip_29_16,ip_29_17,ip_29_18,ip_29_19,ip_29_20,ip_29_21,ip_29_22,ip_29_23,ip_29_24,ip_29_25,ip_29_26,ip_29_27,ip_29_28,ip_29_29,ip_29_30,ip_29_31,ip_29_32,ip_29_33,ip_29_34,ip_29_35,ip_29_36,ip_29_37,ip_29_38,ip_29_39,ip_29_40,ip_29_41,ip_29_42,ip_29_43,ip_29_44,ip_29_45,ip_29_46,ip_29_47,ip_29_48,ip_29_49,ip_29_50,ip_29_51,ip_29_52,ip_29_53,ip_29_54,ip_29_55,ip_29_56,ip_29_57,ip_29_58,ip_29_59,ip_29_60,ip_29_61,ip_29_62,ip_29_63,ip_30_0,ip_30_1,ip_30_2,ip_30_3,ip_30_4,ip_30_5,ip_30_6,ip_30_7,ip_30_8,ip_30_9,ip_30_10,ip_30_11,ip_30_12,ip_30_13,ip_30_14,ip_30_15,ip_30_16,ip_30_17,ip_30_18,ip_30_19,ip_30_20,ip_30_21,ip_30_22,ip_30_23,ip_30_24,ip_30_25,ip_30_26,ip_30_27,ip_30_28,ip_30_29,ip_30_30,ip_30_31,ip_30_32,ip_30_33,ip_30_34,ip_30_35,ip_30_36,ip_30_37,ip_30_38,ip_30_39,ip_30_40,ip_30_41,ip_30_42,ip_30_43,ip_30_44,ip_30_45,ip_30_46,ip_30_47,ip_30_48,ip_30_49,ip_30_50,ip_30_51,ip_30_52,ip_30_53,ip_30_54,ip_30_55,ip_30_56,ip_30_57,ip_30_58,ip_30_59,ip_30_60,ip_30_61,ip_30_62,ip_30_63,ip_31_0,ip_31_1,ip_31_2,ip_31_3,ip_31_4,ip_31_5,ip_31_6,ip_31_7,ip_31_8,ip_31_9,ip_31_10,ip_31_11,ip_31_12,ip_31_13,ip_31_14,ip_31_15,ip_31_16,ip_31_17,ip_31_18,ip_31_19,ip_31_20,ip_31_21,ip_31_22,ip_31_23,ip_31_24,ip_31_25,ip_31_26,ip_31_27,ip_31_28,ip_31_29,ip_31_30,ip_31_31,ip_31_32,ip_31_33,ip_31_34,ip_31_35,ip_31_36,ip_31_37,ip_31_38,ip_31_39,ip_31_40,ip_31_41,ip_31_42,ip_31_43,ip_31_44,ip_31_45,ip_31_46,ip_31_47,ip_31_48,ip_31_49,ip_31_50,ip_31_51,ip_31_52,ip_31_53,ip_31_54,ip_31_55,ip_31_56,ip_31_57,ip_31_58,ip_31_59,ip_31_60,ip_31_61,ip_31_62,ip_31_63,ip_32_0,ip_32_1,ip_32_2,ip_32_3,ip_32_4,ip_32_5,ip_32_6,ip_32_7,ip_32_8,ip_32_9,ip_32_10,ip_32_11,ip_32_12,ip_32_13,ip_32_14,ip_32_15,ip_32_16,ip_32_17,ip_32_18,ip_32_19,ip_32_20,ip_32_21,ip_32_22,ip_32_23,ip_32_24,ip_32_25,ip_32_26,ip_32_27,ip_32_28,ip_32_29,ip_32_30,ip_32_31,ip_32_32,ip_32_33,ip_32_34,ip_32_35,ip_32_36,ip_32_37,ip_32_38,ip_32_39,ip_32_40,ip_32_41,ip_32_42,ip_32_43,ip_32_44,ip_32_45,ip_32_46,ip_32_47,ip_32_48,ip_32_49,ip_32_50,ip_32_51,ip_32_52,ip_32_53,ip_32_54,ip_32_55,ip_32_56,ip_32_57,ip_32_58,ip_32_59,ip_32_60,ip_32_61,ip_32_62,ip_32_63,ip_33_0,ip_33_1,ip_33_2,ip_33_3,ip_33_4,ip_33_5,ip_33_6,ip_33_7,ip_33_8,ip_33_9,ip_33_10,ip_33_11,ip_33_12,ip_33_13,ip_33_14,ip_33_15,ip_33_16,ip_33_17,ip_33_18,ip_33_19,ip_33_20,ip_33_21,ip_33_22,ip_33_23,ip_33_24,ip_33_25,ip_33_26,ip_33_27,ip_33_28,ip_33_29,ip_33_30,ip_33_31,ip_33_32,ip_33_33,ip_33_34,ip_33_35,ip_33_36,ip_33_37,ip_33_38,ip_33_39,ip_33_40,ip_33_41,ip_33_42,ip_33_43,ip_33_44,ip_33_45,ip_33_46,ip_33_47,ip_33_48,ip_33_49,ip_33_50,ip_33_51,ip_33_52,ip_33_53,ip_33_54,ip_33_55,ip_33_56,ip_33_57,ip_33_58,ip_33_59,ip_33_60,ip_33_61,ip_33_62,ip_33_63,ip_34_0,ip_34_1,ip_34_2,ip_34_3,ip_34_4,ip_34_5,ip_34_6,ip_34_7,ip_34_8,ip_34_9,ip_34_10,ip_34_11,ip_34_12,ip_34_13,ip_34_14,ip_34_15,ip_34_16,ip_34_17,ip_34_18,ip_34_19,ip_34_20,ip_34_21,ip_34_22,ip_34_23,ip_34_24,ip_34_25,ip_34_26,ip_34_27,ip_34_28,ip_34_29,ip_34_30,ip_34_31,ip_34_32,ip_34_33,ip_34_34,ip_34_35,ip_34_36,ip_34_37,ip_34_38,ip_34_39,ip_34_40,ip_34_41,ip_34_42,ip_34_43,ip_34_44,ip_34_45,ip_34_46,ip_34_47,ip_34_48,ip_34_49,ip_34_50,ip_34_51,ip_34_52,ip_34_53,ip_34_54,ip_34_55,ip_34_56,ip_34_57,ip_34_58,ip_34_59,ip_34_60,ip_34_61,ip_34_62,ip_34_63,ip_35_0,ip_35_1,ip_35_2,ip_35_3,ip_35_4,ip_35_5,ip_35_6,ip_35_7,ip_35_8,ip_35_9,ip_35_10,ip_35_11,ip_35_12,ip_35_13,ip_35_14,ip_35_15,ip_35_16,ip_35_17,ip_35_18,ip_35_19,ip_35_20,ip_35_21,ip_35_22,ip_35_23,ip_35_24,ip_35_25,ip_35_26,ip_35_27,ip_35_28,ip_35_29,ip_35_30,ip_35_31,ip_35_32,ip_35_33,ip_35_34,ip_35_35,ip_35_36,ip_35_37,ip_35_38,ip_35_39,ip_35_40,ip_35_41,ip_35_42,ip_35_43,ip_35_44,ip_35_45,ip_35_46,ip_35_47,ip_35_48,ip_35_49,ip_35_50,ip_35_51,ip_35_52,ip_35_53,ip_35_54,ip_35_55,ip_35_56,ip_35_57,ip_35_58,ip_35_59,ip_35_60,ip_35_61,ip_35_62,ip_35_63,ip_36_0,ip_36_1,ip_36_2,ip_36_3,ip_36_4,ip_36_5,ip_36_6,ip_36_7,ip_36_8,ip_36_9,ip_36_10,ip_36_11,ip_36_12,ip_36_13,ip_36_14,ip_36_15,ip_36_16,ip_36_17,ip_36_18,ip_36_19,ip_36_20,ip_36_21,ip_36_22,ip_36_23,ip_36_24,ip_36_25,ip_36_26,ip_36_27,ip_36_28,ip_36_29,ip_36_30,ip_36_31,ip_36_32,ip_36_33,ip_36_34,ip_36_35,ip_36_36,ip_36_37,ip_36_38,ip_36_39,ip_36_40,ip_36_41,ip_36_42,ip_36_43,ip_36_44,ip_36_45,ip_36_46,ip_36_47,ip_36_48,ip_36_49,ip_36_50,ip_36_51,ip_36_52,ip_36_53,ip_36_54,ip_36_55,ip_36_56,ip_36_57,ip_36_58,ip_36_59,ip_36_60,ip_36_61,ip_36_62,ip_36_63,ip_37_0,ip_37_1,ip_37_2,ip_37_3,ip_37_4,ip_37_5,ip_37_6,ip_37_7,ip_37_8,ip_37_9,ip_37_10,ip_37_11,ip_37_12,ip_37_13,ip_37_14,ip_37_15,ip_37_16,ip_37_17,ip_37_18,ip_37_19,ip_37_20,ip_37_21,ip_37_22,ip_37_23,ip_37_24,ip_37_25,ip_37_26,ip_37_27,ip_37_28,ip_37_29,ip_37_30,ip_37_31,ip_37_32,ip_37_33,ip_37_34,ip_37_35,ip_37_36,ip_37_37,ip_37_38,ip_37_39,ip_37_40,ip_37_41,ip_37_42,ip_37_43,ip_37_44,ip_37_45,ip_37_46,ip_37_47,ip_37_48,ip_37_49,ip_37_50,ip_37_51,ip_37_52,ip_37_53,ip_37_54,ip_37_55,ip_37_56,ip_37_57,ip_37_58,ip_37_59,ip_37_60,ip_37_61,ip_37_62,ip_37_63,ip_38_0,ip_38_1,ip_38_2,ip_38_3,ip_38_4,ip_38_5,ip_38_6,ip_38_7,ip_38_8,ip_38_9,ip_38_10,ip_38_11,ip_38_12,ip_38_13,ip_38_14,ip_38_15,ip_38_16,ip_38_17,ip_38_18,ip_38_19,ip_38_20,ip_38_21,ip_38_22,ip_38_23,ip_38_24,ip_38_25,ip_38_26,ip_38_27,ip_38_28,ip_38_29,ip_38_30,ip_38_31,ip_38_32,ip_38_33,ip_38_34,ip_38_35,ip_38_36,ip_38_37,ip_38_38,ip_38_39,ip_38_40,ip_38_41,ip_38_42,ip_38_43,ip_38_44,ip_38_45,ip_38_46,ip_38_47,ip_38_48,ip_38_49,ip_38_50,ip_38_51,ip_38_52,ip_38_53,ip_38_54,ip_38_55,ip_38_56,ip_38_57,ip_38_58,ip_38_59,ip_38_60,ip_38_61,ip_38_62,ip_38_63,ip_39_0,ip_39_1,ip_39_2,ip_39_3,ip_39_4,ip_39_5,ip_39_6,ip_39_7,ip_39_8,ip_39_9,ip_39_10,ip_39_11,ip_39_12,ip_39_13,ip_39_14,ip_39_15,ip_39_16,ip_39_17,ip_39_18,ip_39_19,ip_39_20,ip_39_21,ip_39_22,ip_39_23,ip_39_24,ip_39_25,ip_39_26,ip_39_27,ip_39_28,ip_39_29,ip_39_30,ip_39_31,ip_39_32,ip_39_33,ip_39_34,ip_39_35,ip_39_36,ip_39_37,ip_39_38,ip_39_39,ip_39_40,ip_39_41,ip_39_42,ip_39_43,ip_39_44,ip_39_45,ip_39_46,ip_39_47,ip_39_48,ip_39_49,ip_39_50,ip_39_51,ip_39_52,ip_39_53,ip_39_54,ip_39_55,ip_39_56,ip_39_57,ip_39_58,ip_39_59,ip_39_60,ip_39_61,ip_39_62,ip_39_63,ip_40_0,ip_40_1,ip_40_2,ip_40_3,ip_40_4,ip_40_5,ip_40_6,ip_40_7,ip_40_8,ip_40_9,ip_40_10,ip_40_11,ip_40_12,ip_40_13,ip_40_14,ip_40_15,ip_40_16,ip_40_17,ip_40_18,ip_40_19,ip_40_20,ip_40_21,ip_40_22,ip_40_23,ip_40_24,ip_40_25,ip_40_26,ip_40_27,ip_40_28,ip_40_29,ip_40_30,ip_40_31,ip_40_32,ip_40_33,ip_40_34,ip_40_35,ip_40_36,ip_40_37,ip_40_38,ip_40_39,ip_40_40,ip_40_41,ip_40_42,ip_40_43,ip_40_44,ip_40_45,ip_40_46,ip_40_47,ip_40_48,ip_40_49,ip_40_50,ip_40_51,ip_40_52,ip_40_53,ip_40_54,ip_40_55,ip_40_56,ip_40_57,ip_40_58,ip_40_59,ip_40_60,ip_40_61,ip_40_62,ip_40_63,ip_41_0,ip_41_1,ip_41_2,ip_41_3,ip_41_4,ip_41_5,ip_41_6,ip_41_7,ip_41_8,ip_41_9,ip_41_10,ip_41_11,ip_41_12,ip_41_13,ip_41_14,ip_41_15,ip_41_16,ip_41_17,ip_41_18,ip_41_19,ip_41_20,ip_41_21,ip_41_22,ip_41_23,ip_41_24,ip_41_25,ip_41_26,ip_41_27,ip_41_28,ip_41_29,ip_41_30,ip_41_31,ip_41_32,ip_41_33,ip_41_34,ip_41_35,ip_41_36,ip_41_37,ip_41_38,ip_41_39,ip_41_40,ip_41_41,ip_41_42,ip_41_43,ip_41_44,ip_41_45,ip_41_46,ip_41_47,ip_41_48,ip_41_49,ip_41_50,ip_41_51,ip_41_52,ip_41_53,ip_41_54,ip_41_55,ip_41_56,ip_41_57,ip_41_58,ip_41_59,ip_41_60,ip_41_61,ip_41_62,ip_41_63,ip_42_0,ip_42_1,ip_42_2,ip_42_3,ip_42_4,ip_42_5,ip_42_6,ip_42_7,ip_42_8,ip_42_9,ip_42_10,ip_42_11,ip_42_12,ip_42_13,ip_42_14,ip_42_15,ip_42_16,ip_42_17,ip_42_18,ip_42_19,ip_42_20,ip_42_21,ip_42_22,ip_42_23,ip_42_24,ip_42_25,ip_42_26,ip_42_27,ip_42_28,ip_42_29,ip_42_30,ip_42_31,ip_42_32,ip_42_33,ip_42_34,ip_42_35,ip_42_36,ip_42_37,ip_42_38,ip_42_39,ip_42_40,ip_42_41,ip_42_42,ip_42_43,ip_42_44,ip_42_45,ip_42_46,ip_42_47,ip_42_48,ip_42_49,ip_42_50,ip_42_51,ip_42_52,ip_42_53,ip_42_54,ip_42_55,ip_42_56,ip_42_57,ip_42_58,ip_42_59,ip_42_60,ip_42_61,ip_42_62,ip_42_63,ip_43_0,ip_43_1,ip_43_2,ip_43_3,ip_43_4,ip_43_5,ip_43_6,ip_43_7,ip_43_8,ip_43_9,ip_43_10,ip_43_11,ip_43_12,ip_43_13,ip_43_14,ip_43_15,ip_43_16,ip_43_17,ip_43_18,ip_43_19,ip_43_20,ip_43_21,ip_43_22,ip_43_23,ip_43_24,ip_43_25,ip_43_26,ip_43_27,ip_43_28,ip_43_29,ip_43_30,ip_43_31,ip_43_32,ip_43_33,ip_43_34,ip_43_35,ip_43_36,ip_43_37,ip_43_38,ip_43_39,ip_43_40,ip_43_41,ip_43_42,ip_43_43,ip_43_44,ip_43_45,ip_43_46,ip_43_47,ip_43_48,ip_43_49,ip_43_50,ip_43_51,ip_43_52,ip_43_53,ip_43_54,ip_43_55,ip_43_56,ip_43_57,ip_43_58,ip_43_59,ip_43_60,ip_43_61,ip_43_62,ip_43_63,ip_44_0,ip_44_1,ip_44_2,ip_44_3,ip_44_4,ip_44_5,ip_44_6,ip_44_7,ip_44_8,ip_44_9,ip_44_10,ip_44_11,ip_44_12,ip_44_13,ip_44_14,ip_44_15,ip_44_16,ip_44_17,ip_44_18,ip_44_19,ip_44_20,ip_44_21,ip_44_22,ip_44_23,ip_44_24,ip_44_25,ip_44_26,ip_44_27,ip_44_28,ip_44_29,ip_44_30,ip_44_31,ip_44_32,ip_44_33,ip_44_34,ip_44_35,ip_44_36,ip_44_37,ip_44_38,ip_44_39,ip_44_40,ip_44_41,ip_44_42,ip_44_43,ip_44_44,ip_44_45,ip_44_46,ip_44_47,ip_44_48,ip_44_49,ip_44_50,ip_44_51,ip_44_52,ip_44_53,ip_44_54,ip_44_55,ip_44_56,ip_44_57,ip_44_58,ip_44_59,ip_44_60,ip_44_61,ip_44_62,ip_44_63,ip_45_0,ip_45_1,ip_45_2,ip_45_3,ip_45_4,ip_45_5,ip_45_6,ip_45_7,ip_45_8,ip_45_9,ip_45_10,ip_45_11,ip_45_12,ip_45_13,ip_45_14,ip_45_15,ip_45_16,ip_45_17,ip_45_18,ip_45_19,ip_45_20,ip_45_21,ip_45_22,ip_45_23,ip_45_24,ip_45_25,ip_45_26,ip_45_27,ip_45_28,ip_45_29,ip_45_30,ip_45_31,ip_45_32,ip_45_33,ip_45_34,ip_45_35,ip_45_36,ip_45_37,ip_45_38,ip_45_39,ip_45_40,ip_45_41,ip_45_42,ip_45_43,ip_45_44,ip_45_45,ip_45_46,ip_45_47,ip_45_48,ip_45_49,ip_45_50,ip_45_51,ip_45_52,ip_45_53,ip_45_54,ip_45_55,ip_45_56,ip_45_57,ip_45_58,ip_45_59,ip_45_60,ip_45_61,ip_45_62,ip_45_63,ip_46_0,ip_46_1,ip_46_2,ip_46_3,ip_46_4,ip_46_5,ip_46_6,ip_46_7,ip_46_8,ip_46_9,ip_46_10,ip_46_11,ip_46_12,ip_46_13,ip_46_14,ip_46_15,ip_46_16,ip_46_17,ip_46_18,ip_46_19,ip_46_20,ip_46_21,ip_46_22,ip_46_23,ip_46_24,ip_46_25,ip_46_26,ip_46_27,ip_46_28,ip_46_29,ip_46_30,ip_46_31,ip_46_32,ip_46_33,ip_46_34,ip_46_35,ip_46_36,ip_46_37,ip_46_38,ip_46_39,ip_46_40,ip_46_41,ip_46_42,ip_46_43,ip_46_44,ip_46_45,ip_46_46,ip_46_47,ip_46_48,ip_46_49,ip_46_50,ip_46_51,ip_46_52,ip_46_53,ip_46_54,ip_46_55,ip_46_56,ip_46_57,ip_46_58,ip_46_59,ip_46_60,ip_46_61,ip_46_62,ip_46_63,ip_47_0,ip_47_1,ip_47_2,ip_47_3,ip_47_4,ip_47_5,ip_47_6,ip_47_7,ip_47_8,ip_47_9,ip_47_10,ip_47_11,ip_47_12,ip_47_13,ip_47_14,ip_47_15,ip_47_16,ip_47_17,ip_47_18,ip_47_19,ip_47_20,ip_47_21,ip_47_22,ip_47_23,ip_47_24,ip_47_25,ip_47_26,ip_47_27,ip_47_28,ip_47_29,ip_47_30,ip_47_31,ip_47_32,ip_47_33,ip_47_34,ip_47_35,ip_47_36,ip_47_37,ip_47_38,ip_47_39,ip_47_40,ip_47_41,ip_47_42,ip_47_43,ip_47_44,ip_47_45,ip_47_46,ip_47_47,ip_47_48,ip_47_49,ip_47_50,ip_47_51,ip_47_52,ip_47_53,ip_47_54,ip_47_55,ip_47_56,ip_47_57,ip_47_58,ip_47_59,ip_47_60,ip_47_61,ip_47_62,ip_47_63,ip_48_0,ip_48_1,ip_48_2,ip_48_3,ip_48_4,ip_48_5,ip_48_6,ip_48_7,ip_48_8,ip_48_9,ip_48_10,ip_48_11,ip_48_12,ip_48_13,ip_48_14,ip_48_15,ip_48_16,ip_48_17,ip_48_18,ip_48_19,ip_48_20,ip_48_21,ip_48_22,ip_48_23,ip_48_24,ip_48_25,ip_48_26,ip_48_27,ip_48_28,ip_48_29,ip_48_30,ip_48_31,ip_48_32,ip_48_33,ip_48_34,ip_48_35,ip_48_36,ip_48_37,ip_48_38,ip_48_39,ip_48_40,ip_48_41,ip_48_42,ip_48_43,ip_48_44,ip_48_45,ip_48_46,ip_48_47,ip_48_48,ip_48_49,ip_48_50,ip_48_51,ip_48_52,ip_48_53,ip_48_54,ip_48_55,ip_48_56,ip_48_57,ip_48_58,ip_48_59,ip_48_60,ip_48_61,ip_48_62,ip_48_63,ip_49_0,ip_49_1,ip_49_2,ip_49_3,ip_49_4,ip_49_5,ip_49_6,ip_49_7,ip_49_8,ip_49_9,ip_49_10,ip_49_11,ip_49_12,ip_49_13,ip_49_14,ip_49_15,ip_49_16,ip_49_17,ip_49_18,ip_49_19,ip_49_20,ip_49_21,ip_49_22,ip_49_23,ip_49_24,ip_49_25,ip_49_26,ip_49_27,ip_49_28,ip_49_29,ip_49_30,ip_49_31,ip_49_32,ip_49_33,ip_49_34,ip_49_35,ip_49_36,ip_49_37,ip_49_38,ip_49_39,ip_49_40,ip_49_41,ip_49_42,ip_49_43,ip_49_44,ip_49_45,ip_49_46,ip_49_47,ip_49_48,ip_49_49,ip_49_50,ip_49_51,ip_49_52,ip_49_53,ip_49_54,ip_49_55,ip_49_56,ip_49_57,ip_49_58,ip_49_59,ip_49_60,ip_49_61,ip_49_62,ip_49_63,ip_50_0,ip_50_1,ip_50_2,ip_50_3,ip_50_4,ip_50_5,ip_50_6,ip_50_7,ip_50_8,ip_50_9,ip_50_10,ip_50_11,ip_50_12,ip_50_13,ip_50_14,ip_50_15,ip_50_16,ip_50_17,ip_50_18,ip_50_19,ip_50_20,ip_50_21,ip_50_22,ip_50_23,ip_50_24,ip_50_25,ip_50_26,ip_50_27,ip_50_28,ip_50_29,ip_50_30,ip_50_31,ip_50_32,ip_50_33,ip_50_34,ip_50_35,ip_50_36,ip_50_37,ip_50_38,ip_50_39,ip_50_40,ip_50_41,ip_50_42,ip_50_43,ip_50_44,ip_50_45,ip_50_46,ip_50_47,ip_50_48,ip_50_49,ip_50_50,ip_50_51,ip_50_52,ip_50_53,ip_50_54,ip_50_55,ip_50_56,ip_50_57,ip_50_58,ip_50_59,ip_50_60,ip_50_61,ip_50_62,ip_50_63,ip_51_0,ip_51_1,ip_51_2,ip_51_3,ip_51_4,ip_51_5,ip_51_6,ip_51_7,ip_51_8,ip_51_9,ip_51_10,ip_51_11,ip_51_12,ip_51_13,ip_51_14,ip_51_15,ip_51_16,ip_51_17,ip_51_18,ip_51_19,ip_51_20,ip_51_21,ip_51_22,ip_51_23,ip_51_24,ip_51_25,ip_51_26,ip_51_27,ip_51_28,ip_51_29,ip_51_30,ip_51_31,ip_51_32,ip_51_33,ip_51_34,ip_51_35,ip_51_36,ip_51_37,ip_51_38,ip_51_39,ip_51_40,ip_51_41,ip_51_42,ip_51_43,ip_51_44,ip_51_45,ip_51_46,ip_51_47,ip_51_48,ip_51_49,ip_51_50,ip_51_51,ip_51_52,ip_51_53,ip_51_54,ip_51_55,ip_51_56,ip_51_57,ip_51_58,ip_51_59,ip_51_60,ip_51_61,ip_51_62,ip_51_63,ip_52_0,ip_52_1,ip_52_2,ip_52_3,ip_52_4,ip_52_5,ip_52_6,ip_52_7,ip_52_8,ip_52_9,ip_52_10,ip_52_11,ip_52_12,ip_52_13,ip_52_14,ip_52_15,ip_52_16,ip_52_17,ip_52_18,ip_52_19,ip_52_20,ip_52_21,ip_52_22,ip_52_23,ip_52_24,ip_52_25,ip_52_26,ip_52_27,ip_52_28,ip_52_29,ip_52_30,ip_52_31,ip_52_32,ip_52_33,ip_52_34,ip_52_35,ip_52_36,ip_52_37,ip_52_38,ip_52_39,ip_52_40,ip_52_41,ip_52_42,ip_52_43,ip_52_44,ip_52_45,ip_52_46,ip_52_47,ip_52_48,ip_52_49,ip_52_50,ip_52_51,ip_52_52,ip_52_53,ip_52_54,ip_52_55,ip_52_56,ip_52_57,ip_52_58,ip_52_59,ip_52_60,ip_52_61,ip_52_62,ip_52_63,ip_53_0,ip_53_1,ip_53_2,ip_53_3,ip_53_4,ip_53_5,ip_53_6,ip_53_7,ip_53_8,ip_53_9,ip_53_10,ip_53_11,ip_53_12,ip_53_13,ip_53_14,ip_53_15,ip_53_16,ip_53_17,ip_53_18,ip_53_19,ip_53_20,ip_53_21,ip_53_22,ip_53_23,ip_53_24,ip_53_25,ip_53_26,ip_53_27,ip_53_28,ip_53_29,ip_53_30,ip_53_31,ip_53_32,ip_53_33,ip_53_34,ip_53_35,ip_53_36,ip_53_37,ip_53_38,ip_53_39,ip_53_40,ip_53_41,ip_53_42,ip_53_43,ip_53_44,ip_53_45,ip_53_46,ip_53_47,ip_53_48,ip_53_49,ip_53_50,ip_53_51,ip_53_52,ip_53_53,ip_53_54,ip_53_55,ip_53_56,ip_53_57,ip_53_58,ip_53_59,ip_53_60,ip_53_61,ip_53_62,ip_53_63,ip_54_0,ip_54_1,ip_54_2,ip_54_3,ip_54_4,ip_54_5,ip_54_6,ip_54_7,ip_54_8,ip_54_9,ip_54_10,ip_54_11,ip_54_12,ip_54_13,ip_54_14,ip_54_15,ip_54_16,ip_54_17,ip_54_18,ip_54_19,ip_54_20,ip_54_21,ip_54_22,ip_54_23,ip_54_24,ip_54_25,ip_54_26,ip_54_27,ip_54_28,ip_54_29,ip_54_30,ip_54_31,ip_54_32,ip_54_33,ip_54_34,ip_54_35,ip_54_36,ip_54_37,ip_54_38,ip_54_39,ip_54_40,ip_54_41,ip_54_42,ip_54_43,ip_54_44,ip_54_45,ip_54_46,ip_54_47,ip_54_48,ip_54_49,ip_54_50,ip_54_51,ip_54_52,ip_54_53,ip_54_54,ip_54_55,ip_54_56,ip_54_57,ip_54_58,ip_54_59,ip_54_60,ip_54_61,ip_54_62,ip_54_63,ip_55_0,ip_55_1,ip_55_2,ip_55_3,ip_55_4,ip_55_5,ip_55_6,ip_55_7,ip_55_8,ip_55_9,ip_55_10,ip_55_11,ip_55_12,ip_55_13,ip_55_14,ip_55_15,ip_55_16,ip_55_17,ip_55_18,ip_55_19,ip_55_20,ip_55_21,ip_55_22,ip_55_23,ip_55_24,ip_55_25,ip_55_26,ip_55_27,ip_55_28,ip_55_29,ip_55_30,ip_55_31,ip_55_32,ip_55_33,ip_55_34,ip_55_35,ip_55_36,ip_55_37,ip_55_38,ip_55_39,ip_55_40,ip_55_41,ip_55_42,ip_55_43,ip_55_44,ip_55_45,ip_55_46,ip_55_47,ip_55_48,ip_55_49,ip_55_50,ip_55_51,ip_55_52,ip_55_53,ip_55_54,ip_55_55,ip_55_56,ip_55_57,ip_55_58,ip_55_59,ip_55_60,ip_55_61,ip_55_62,ip_55_63,ip_56_0,ip_56_1,ip_56_2,ip_56_3,ip_56_4,ip_56_5,ip_56_6,ip_56_7,ip_56_8,ip_56_9,ip_56_10,ip_56_11,ip_56_12,ip_56_13,ip_56_14,ip_56_15,ip_56_16,ip_56_17,ip_56_18,ip_56_19,ip_56_20,ip_56_21,ip_56_22,ip_56_23,ip_56_24,ip_56_25,ip_56_26,ip_56_27,ip_56_28,ip_56_29,ip_56_30,ip_56_31,ip_56_32,ip_56_33,ip_56_34,ip_56_35,ip_56_36,ip_56_37,ip_56_38,ip_56_39,ip_56_40,ip_56_41,ip_56_42,ip_56_43,ip_56_44,ip_56_45,ip_56_46,ip_56_47,ip_56_48,ip_56_49,ip_56_50,ip_56_51,ip_56_52,ip_56_53,ip_56_54,ip_56_55,ip_56_56,ip_56_57,ip_56_58,ip_56_59,ip_56_60,ip_56_61,ip_56_62,ip_56_63,ip_57_0,ip_57_1,ip_57_2,ip_57_3,ip_57_4,ip_57_5,ip_57_6,ip_57_7,ip_57_8,ip_57_9,ip_57_10,ip_57_11,ip_57_12,ip_57_13,ip_57_14,ip_57_15,ip_57_16,ip_57_17,ip_57_18,ip_57_19,ip_57_20,ip_57_21,ip_57_22,ip_57_23,ip_57_24,ip_57_25,ip_57_26,ip_57_27,ip_57_28,ip_57_29,ip_57_30,ip_57_31,ip_57_32,ip_57_33,ip_57_34,ip_57_35,ip_57_36,ip_57_37,ip_57_38,ip_57_39,ip_57_40,ip_57_41,ip_57_42,ip_57_43,ip_57_44,ip_57_45,ip_57_46,ip_57_47,ip_57_48,ip_57_49,ip_57_50,ip_57_51,ip_57_52,ip_57_53,ip_57_54,ip_57_55,ip_57_56,ip_57_57,ip_57_58,ip_57_59,ip_57_60,ip_57_61,ip_57_62,ip_57_63,ip_58_0,ip_58_1,ip_58_2,ip_58_3,ip_58_4,ip_58_5,ip_58_6,ip_58_7,ip_58_8,ip_58_9,ip_58_10,ip_58_11,ip_58_12,ip_58_13,ip_58_14,ip_58_15,ip_58_16,ip_58_17,ip_58_18,ip_58_19,ip_58_20,ip_58_21,ip_58_22,ip_58_23,ip_58_24,ip_58_25,ip_58_26,ip_58_27,ip_58_28,ip_58_29,ip_58_30,ip_58_31,ip_58_32,ip_58_33,ip_58_34,ip_58_35,ip_58_36,ip_58_37,ip_58_38,ip_58_39,ip_58_40,ip_58_41,ip_58_42,ip_58_43,ip_58_44,ip_58_45,ip_58_46,ip_58_47,ip_58_48,ip_58_49,ip_58_50,ip_58_51,ip_58_52,ip_58_53,ip_58_54,ip_58_55,ip_58_56,ip_58_57,ip_58_58,ip_58_59,ip_58_60,ip_58_61,ip_58_62,ip_58_63,ip_59_0,ip_59_1,ip_59_2,ip_59_3,ip_59_4,ip_59_5,ip_59_6,ip_59_7,ip_59_8,ip_59_9,ip_59_10,ip_59_11,ip_59_12,ip_59_13,ip_59_14,ip_59_15,ip_59_16,ip_59_17,ip_59_18,ip_59_19,ip_59_20,ip_59_21,ip_59_22,ip_59_23,ip_59_24,ip_59_25,ip_59_26,ip_59_27,ip_59_28,ip_59_29,ip_59_30,ip_59_31,ip_59_32,ip_59_33,ip_59_34,ip_59_35,ip_59_36,ip_59_37,ip_59_38,ip_59_39,ip_59_40,ip_59_41,ip_59_42,ip_59_43,ip_59_44,ip_59_45,ip_59_46,ip_59_47,ip_59_48,ip_59_49,ip_59_50,ip_59_51,ip_59_52,ip_59_53,ip_59_54,ip_59_55,ip_59_56,ip_59_57,ip_59_58,ip_59_59,ip_59_60,ip_59_61,ip_59_62,ip_59_63,ip_60_0,ip_60_1,ip_60_2,ip_60_3,ip_60_4,ip_60_5,ip_60_6,ip_60_7,ip_60_8,ip_60_9,ip_60_10,ip_60_11,ip_60_12,ip_60_13,ip_60_14,ip_60_15,ip_60_16,ip_60_17,ip_60_18,ip_60_19,ip_60_20,ip_60_21,ip_60_22,ip_60_23,ip_60_24,ip_60_25,ip_60_26,ip_60_27,ip_60_28,ip_60_29,ip_60_30,ip_60_31,ip_60_32,ip_60_33,ip_60_34,ip_60_35,ip_60_36,ip_60_37,ip_60_38,ip_60_39,ip_60_40,ip_60_41,ip_60_42,ip_60_43,ip_60_44,ip_60_45,ip_60_46,ip_60_47,ip_60_48,ip_60_49,ip_60_50,ip_60_51,ip_60_52,ip_60_53,ip_60_54,ip_60_55,ip_60_56,ip_60_57,ip_60_58,ip_60_59,ip_60_60,ip_60_61,ip_60_62,ip_60_63,ip_61_0,ip_61_1,ip_61_2,ip_61_3,ip_61_4,ip_61_5,ip_61_6,ip_61_7,ip_61_8,ip_61_9,ip_61_10,ip_61_11,ip_61_12,ip_61_13,ip_61_14,ip_61_15,ip_61_16,ip_61_17,ip_61_18,ip_61_19,ip_61_20,ip_61_21,ip_61_22,ip_61_23,ip_61_24,ip_61_25,ip_61_26,ip_61_27,ip_61_28,ip_61_29,ip_61_30,ip_61_31,ip_61_32,ip_61_33,ip_61_34,ip_61_35,ip_61_36,ip_61_37,ip_61_38,ip_61_39,ip_61_40,ip_61_41,ip_61_42,ip_61_43,ip_61_44,ip_61_45,ip_61_46,ip_61_47,ip_61_48,ip_61_49,ip_61_50,ip_61_51,ip_61_52,ip_61_53,ip_61_54,ip_61_55,ip_61_56,ip_61_57,ip_61_58,ip_61_59,ip_61_60,ip_61_61,ip_61_62,ip_61_63,ip_62_0,ip_62_1,ip_62_2,ip_62_3,ip_62_4,ip_62_5,ip_62_6,ip_62_7,ip_62_8,ip_62_9,ip_62_10,ip_62_11,ip_62_12,ip_62_13,ip_62_14,ip_62_15,ip_62_16,ip_62_17,ip_62_18,ip_62_19,ip_62_20,ip_62_21,ip_62_22,ip_62_23,ip_62_24,ip_62_25,ip_62_26,ip_62_27,ip_62_28,ip_62_29,ip_62_30,ip_62_31,ip_62_32,ip_62_33,ip_62_34,ip_62_35,ip_62_36,ip_62_37,ip_62_38,ip_62_39,ip_62_40,ip_62_41,ip_62_42,ip_62_43,ip_62_44,ip_62_45,ip_62_46,ip_62_47,ip_62_48,ip_62_49,ip_62_50,ip_62_51,ip_62_52,ip_62_53,ip_62_54,ip_62_55,ip_62_56,ip_62_57,ip_62_58,ip_62_59,ip_62_60,ip_62_61,ip_62_62,ip_62_63,ip_63_0,ip_63_1,ip_63_2,ip_63_3,ip_63_4,ip_63_5,ip_63_6,ip_63_7,ip_63_8,ip_63_9,ip_63_10,ip_63_11,ip_63_12,ip_63_13,ip_63_14,ip_63_15,ip_63_16,ip_63_17,ip_63_18,ip_63_19,ip_63_20,ip_63_21,ip_63_22,ip_63_23,ip_63_24,ip_63_25,ip_63_26,ip_63_27,ip_63_28,ip_63_29,ip_63_30,ip_63_31,ip_63_32,ip_63_33,ip_63_34,ip_63_35,ip_63_36,ip_63_37,ip_63_38,ip_63_39,ip_63_40,ip_63_41,ip_63_42,ip_63_43,ip_63_44,ip_63_45,ip_63_46,ip_63_47,ip_63_48,ip_63_49,ip_63_50,ip_63_51,ip_63_52,ip_63_53,ip_63_54,ip_63_55,ip_63_56,ip_63_57,ip_63_58,ip_63_59,ip_63_60,ip_63_61,ip_63_62,ip_63_63;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149,p1150,p1151,p1152,p1153,p1154,p1155,p1156,p1157,p1158,p1159,p1160,p1161,p1162,p1163,p1164,p1165,p1166,p1167,p1168,p1169,p1170,p1171,p1172,p1173,p1174,p1175,p1176,p1177,p1178,p1179,p1180,p1181,p1182,p1183,p1184,p1185,p1186,p1187,p1188,p1189,p1190,p1191,p1192,p1193,p1194,p1195,p1196,p1197,p1198,p1199,p1200,p1201,p1202,p1203,p1204,p1205,p1206,p1207,p1208,p1209,p1210,p1211,p1212,p1213,p1214,p1215,p1216,p1217,p1218,p1219,p1220,p1221,p1222,p1223,p1224,p1225,p1226,p1227,p1228,p1229,p1230,p1231,p1232,p1233,p1234,p1235,p1236,p1237,p1238,p1239,p1240,p1241,p1242,p1243,p1244,p1245,p1246,p1247,p1248,p1249,p1250,p1251,p1252,p1253,p1254,p1255,p1256,p1257,p1258,p1259,p1260,p1261,p1262,p1263,p1264,p1265,p1266,p1267,p1268,p1269,p1270,p1271,p1272,p1273,p1274,p1275,p1276,p1277,p1278,p1279,p1280,p1281,p1282,p1283,p1284,p1285,p1286,p1287,p1288,p1289,p1290,p1291,p1292,p1293,p1294,p1295,p1296,p1297,p1298,p1299,p1300,p1301,p1302,p1303,p1304,p1305,p1306,p1307,p1308,p1309,p1310,p1311,p1312,p1313,p1314,p1315,p1316,p1317,p1318,p1319,p1320,p1321,p1322,p1323,p1324,p1325,p1326,p1327,p1328,p1329,p1330,p1331,p1332,p1333,p1334,p1335,p1336,p1337,p1338,p1339,p1340,p1341,p1342,p1343,p1344,p1345,p1346,p1347,p1348,p1349,p1350,p1351,p1352,p1353,p1354,p1355,p1356,p1357,p1358,p1359,p1360,p1361,p1362,p1363,p1364,p1365,p1366,p1367,p1368,p1369,p1370,p1371,p1372,p1373,p1374,p1375,p1376,p1377,p1378,p1379,p1380,p1381,p1382,p1383,p1384,p1385,p1386,p1387,p1388,p1389,p1390,p1391,p1392,p1393,p1394,p1395,p1396,p1397,p1398,p1399,p1400,p1401,p1402,p1403,p1404,p1405,p1406,p1407,p1408,p1409,p1410,p1411,p1412,p1413,p1414,p1415,p1416,p1417,p1418,p1419,p1420,p1421,p1422,p1423,p1424,p1425,p1426,p1427,p1428,p1429,p1430,p1431,p1432,p1433,p1434,p1435,p1436,p1437,p1438,p1439,p1440,p1441,p1442,p1443,p1444,p1445,p1446,p1447,p1448,p1449,p1450,p1451,p1452,p1453,p1454,p1455,p1456,p1457,p1458,p1459,p1460,p1461,p1462,p1463,p1464,p1465,p1466,p1467,p1468,p1469,p1470,p1471,p1472,p1473,p1474,p1475,p1476,p1477,p1478,p1479,p1480,p1481,p1482,p1483,p1484,p1485,p1486,p1487,p1488,p1489,p1490,p1491,p1492,p1493,p1494,p1495,p1496,p1497,p1498,p1499,p1500,p1501,p1502,p1503,p1504,p1505,p1506,p1507,p1508,p1509,p1510,p1511,p1512,p1513,p1514,p1515,p1516,p1517,p1518,p1519,p1520,p1521,p1522,p1523,p1524,p1525,p1526,p1527,p1528,p1529,p1530,p1531,p1532,p1533,p1534,p1535,p1536,p1537,p1538,p1539,p1540,p1541,p1542,p1543,p1544,p1545,p1546,p1547,p1548,p1549,p1550,p1551,p1552,p1553,p1554,p1555,p1556,p1557,p1558,p1559,p1560,p1561,p1562,p1563,p1564,p1565,p1566,p1567,p1568,p1569,p1570,p1571,p1572,p1573,p1574,p1575,p1576,p1577,p1578,p1579,p1580,p1581,p1582,p1583,p1584,p1585,p1586,p1587,p1588,p1589,p1590,p1591,p1592,p1593,p1594,p1595,p1596,p1597,p1598,p1599,p1600,p1601,p1602,p1603,p1604,p1605,p1606,p1607,p1608,p1609,p1610,p1611,p1612,p1613,p1614,p1615,p1616,p1617,p1618,p1619,p1620,p1621,p1622,p1623,p1624,p1625,p1626,p1627,p1628,p1629,p1630,p1631,p1632,p1633,p1634,p1635,p1636,p1637,p1638,p1639,p1640,p1641,p1642,p1643,p1644,p1645,p1646,p1647,p1648,p1649,p1650,p1651,p1652,p1653,p1654,p1655,p1656,p1657,p1658,p1659,p1660,p1661,p1662,p1663,p1664,p1665,p1666,p1667,p1668,p1669,p1670,p1671,p1672,p1673,p1674,p1675,p1676,p1677,p1678,p1679,p1680,p1681,p1682,p1683,p1684,p1685,p1686,p1687,p1688,p1689,p1690,p1691,p1692,p1693,p1694,p1695,p1696,p1697,p1698,p1699,p1700,p1701,p1702,p1703,p1704,p1705,p1706,p1707,p1708,p1709,p1710,p1711,p1712,p1713,p1714,p1715,p1716,p1717,p1718,p1719,p1720,p1721,p1722,p1723,p1724,p1725,p1726,p1727,p1728,p1729,p1730,p1731,p1732,p1733,p1734,p1735,p1736,p1737,p1738,p1739,p1740,p1741,p1742,p1743,p1744,p1745,p1746,p1747,p1748,p1749,p1750,p1751,p1752,p1753,p1754,p1755,p1756,p1757,p1758,p1759,p1760,p1761,p1762,p1763,p1764,p1765,p1766,p1767,p1768,p1769,p1770,p1771,p1772,p1773,p1774,p1775,p1776,p1777,p1778,p1779,p1780,p1781,p1782,p1783,p1784,p1785,p1786,p1787,p1788,p1789,p1790,p1791,p1792,p1793,p1794,p1795,p1796,p1797,p1798,p1799,p1800,p1801,p1802,p1803,p1804,p1805,p1806,p1807,p1808,p1809,p1810,p1811,p1812,p1813,p1814,p1815,p1816,p1817,p1818,p1819,p1820,p1821,p1822,p1823,p1824,p1825,p1826,p1827,p1828,p1829,p1830,p1831,p1832,p1833,p1834,p1835,p1836,p1837,p1838,p1839,p1840,p1841,p1842,p1843,p1844,p1845,p1846,p1847,p1848,p1849,p1850,p1851,p1852,p1853,p1854,p1855,p1856,p1857,p1858,p1859,p1860,p1861,p1862,p1863,p1864,p1865,p1866,p1867,p1868,p1869,p1870,p1871,p1872,p1873,p1874,p1875,p1876,p1877,p1878,p1879,p1880,p1881,p1882,p1883,p1884,p1885,p1886,p1887,p1888,p1889,p1890,p1891,p1892,p1893,p1894,p1895,p1896,p1897,p1898,p1899,p1900,p1901,p1902,p1903,p1904,p1905,p1906,p1907,p1908,p1909,p1910,p1911,p1912,p1913,p1914,p1915,p1916,p1917,p1918,p1919,p1920,p1921,p1922,p1923,p1924,p1925,p1926,p1927,p1928,p1929,p1930,p1931,p1932,p1933,p1934,p1935,p1936,p1937,p1938,p1939,p1940,p1941,p1942,p1943,p1944,p1945,p1946,p1947,p1948,p1949,p1950,p1951,p1952,p1953,p1954,p1955,p1956,p1957,p1958,p1959,p1960,p1961,p1962,p1963,p1964,p1965,p1966,p1967,p1968,p1969,p1970,p1971,p1972,p1973,p1974,p1975,p1976,p1977,p1978,p1979,p1980,p1981,p1982,p1983,p1984,p1985,p1986,p1987,p1988,p1989,p1990,p1991,p1992,p1993,p1994,p1995,p1996,p1997,p1998,p1999,p2000,p2001,p2002,p2003,p2004,p2005,p2006,p2007,p2008,p2009,p2010,p2011,p2012,p2013,p2014,p2015,p2016,p2017,p2018,p2019,p2020,p2021,p2022,p2023,p2024,p2025,p2026,p2027,p2028,p2029,p2030,p2031,p2032,p2033,p2034,p2035,p2036,p2037,p2038,p2039,p2040,p2041,p2042,p2043,p2044,p2045,p2046,p2047,p2048,p2049,p2050,p2051,p2052,p2053,p2054,p2055,p2056,p2057,p2058,p2059,p2060,p2061,p2062,p2063,p2064,p2065,p2066,p2067,p2068,p2069,p2070,p2071,p2072,p2073,p2074,p2075,p2076,p2077,p2078,p2079,p2080,p2081,p2082,p2083,p2084,p2085,p2086,p2087,p2088,p2089,p2090,p2091,p2092,p2093,p2094,p2095,p2096,p2097,p2098,p2099,p2100,p2101,p2102,p2103,p2104,p2105,p2106,p2107,p2108,p2109,p2110,p2111,p2112,p2113,p2114,p2115,p2116,p2117,p2118,p2119,p2120,p2121,p2122,p2123,p2124,p2125,p2126,p2127,p2128,p2129,p2130,p2131,p2132,p2133,p2134,p2135,p2136,p2137,p2138,p2139,p2140,p2141,p2142,p2143,p2144,p2145,p2146,p2147,p2148,p2149,p2150,p2151,p2152,p2153,p2154,p2155,p2156,p2157,p2158,p2159,p2160,p2161,p2162,p2163,p2164,p2165,p2166,p2167,p2168,p2169,p2170,p2171,p2172,p2173,p2174,p2175,p2176,p2177,p2178,p2179,p2180,p2181,p2182,p2183,p2184,p2185,p2186,p2187,p2188,p2189,p2190,p2191,p2192,p2193,p2194,p2195,p2196,p2197,p2198,p2199,p2200,p2201,p2202,p2203,p2204,p2205,p2206,p2207,p2208,p2209,p2210,p2211,p2212,p2213,p2214,p2215,p2216,p2217,p2218,p2219,p2220,p2221,p2222,p2223,p2224,p2225,p2226,p2227,p2228,p2229,p2230,p2231,p2232,p2233,p2234,p2235,p2236,p2237,p2238,p2239,p2240,p2241,p2242,p2243,p2244,p2245,p2246,p2247,p2248,p2249,p2250,p2251,p2252,p2253,p2254,p2255,p2256,p2257,p2258,p2259,p2260,p2261,p2262,p2263,p2264,p2265,p2266,p2267,p2268,p2269,p2270,p2271,p2272,p2273,p2274,p2275,p2276,p2277,p2278,p2279,p2280,p2281,p2282,p2283,p2284,p2285,p2286,p2287,p2288,p2289,p2290,p2291,p2292,p2293,p2294,p2295,p2296,p2297,p2298,p2299,p2300,p2301,p2302,p2303,p2304,p2305,p2306,p2307,p2308,p2309,p2310,p2311,p2312,p2313,p2314,p2315,p2316,p2317,p2318,p2319,p2320,p2321,p2322,p2323,p2324,p2325,p2326,p2327,p2328,p2329,p2330,p2331,p2332,p2333,p2334,p2335,p2336,p2337,p2338,p2339,p2340,p2341,p2342,p2343,p2344,p2345,p2346,p2347,p2348,p2349,p2350,p2351,p2352,p2353,p2354,p2355,p2356,p2357,p2358,p2359,p2360,p2361,p2362,p2363,p2364,p2365,p2366,p2367,p2368,p2369,p2370,p2371,p2372,p2373,p2374,p2375,p2376,p2377,p2378,p2379,p2380,p2381,p2382,p2383,p2384,p2385,p2386,p2387,p2388,p2389,p2390,p2391,p2392,p2393,p2394,p2395,p2396,p2397,p2398,p2399,p2400,p2401,p2402,p2403,p2404,p2405,p2406,p2407,p2408,p2409,p2410,p2411,p2412,p2413,p2414,p2415,p2416,p2417,p2418,p2419,p2420,p2421,p2422,p2423,p2424,p2425,p2426,p2427,p2428,p2429,p2430,p2431,p2432,p2433,p2434,p2435,p2436,p2437,p2438,p2439,p2440,p2441,p2442,p2443,p2444,p2445,p2446,p2447,p2448,p2449,p2450,p2451,p2452,p2453,p2454,p2455,p2456,p2457,p2458,p2459,p2460,p2461,p2462,p2463,p2464,p2465,p2466,p2467,p2468,p2469,p2470,p2471,p2472,p2473,p2474,p2475,p2476,p2477,p2478,p2479,p2480,p2481,p2482,p2483,p2484,p2485,p2486,p2487,p2488,p2489,p2490,p2491,p2492,p2493,p2494,p2495,p2496,p2497,p2498,p2499,p2500,p2501,p2502,p2503,p2504,p2505,p2506,p2507,p2508,p2509,p2510,p2511,p2512,p2513,p2514,p2515,p2516,p2517,p2518,p2519,p2520,p2521,p2522,p2523,p2524,p2525,p2526,p2527,p2528,p2529,p2530,p2531,p2532,p2533,p2534,p2535,p2536,p2537,p2538,p2539,p2540,p2541,p2542,p2543,p2544,p2545,p2546,p2547,p2548,p2549,p2550,p2551,p2552,p2553,p2554,p2555,p2556,p2557,p2558,p2559,p2560,p2561,p2562,p2563,p2564,p2565,p2566,p2567,p2568,p2569,p2570,p2571,p2572,p2573,p2574,p2575,p2576,p2577,p2578,p2579,p2580,p2581,p2582,p2583,p2584,p2585,p2586,p2587,p2588,p2589,p2590,p2591,p2592,p2593,p2594,p2595,p2596,p2597,p2598,p2599,p2600,p2601,p2602,p2603,p2604,p2605,p2606,p2607,p2608,p2609,p2610,p2611,p2612,p2613,p2614,p2615,p2616,p2617,p2618,p2619,p2620,p2621,p2622,p2623,p2624,p2625,p2626,p2627,p2628,p2629,p2630,p2631,p2632,p2633,p2634,p2635,p2636,p2637,p2638,p2639,p2640,p2641,p2642,p2643,p2644,p2645,p2646,p2647,p2648,p2649,p2650,p2651,p2652,p2653,p2654,p2655,p2656,p2657,p2658,p2659,p2660,p2661,p2662,p2663,p2664,p2665,p2666,p2667,p2668,p2669,p2670,p2671,p2672,p2673,p2674,p2675,p2676,p2677,p2678,p2679,p2680,p2681,p2682,p2683,p2684,p2685,p2686,p2687,p2688,p2689,p2690,p2691,p2692,p2693,p2694,p2695,p2696,p2697,p2698,p2699,p2700,p2701,p2702,p2703,p2704,p2705,p2706,p2707,p2708,p2709,p2710,p2711,p2712,p2713,p2714,p2715,p2716,p2717,p2718,p2719,p2720,p2721,p2722,p2723,p2724,p2725,p2726,p2727,p2728,p2729,p2730,p2731,p2732,p2733,p2734,p2735,p2736,p2737,p2738,p2739,p2740,p2741,p2742,p2743,p2744,p2745,p2746,p2747,p2748,p2749,p2750,p2751,p2752,p2753,p2754,p2755,p2756,p2757,p2758,p2759,p2760,p2761,p2762,p2763,p2764,p2765,p2766,p2767,p2768,p2769,p2770,p2771,p2772,p2773,p2774,p2775,p2776,p2777,p2778,p2779,p2780,p2781,p2782,p2783,p2784,p2785,p2786,p2787,p2788,p2789,p2790,p2791,p2792,p2793,p2794,p2795,p2796,p2797,p2798,p2799,p2800,p2801,p2802,p2803,p2804,p2805,p2806,p2807,p2808,p2809,p2810,p2811,p2812,p2813,p2814,p2815,p2816,p2817,p2818,p2819,p2820,p2821,p2822,p2823,p2824,p2825,p2826,p2827,p2828,p2829,p2830,p2831,p2832,p2833,p2834,p2835,p2836,p2837,p2838,p2839,p2840,p2841,p2842,p2843,p2844,p2845,p2846,p2847,p2848,p2849,p2850,p2851,p2852,p2853,p2854,p2855,p2856,p2857,p2858,p2859,p2860,p2861,p2862,p2863,p2864,p2865,p2866,p2867,p2868,p2869,p2870,p2871,p2872,p2873,p2874,p2875,p2876,p2877,p2878,p2879,p2880,p2881,p2882,p2883,p2884,p2885,p2886,p2887,p2888,p2889,p2890,p2891,p2892,p2893,p2894,p2895,p2896,p2897,p2898,p2899,p2900,p2901,p2902,p2903,p2904,p2905,p2906,p2907,p2908,p2909,p2910,p2911,p2912,p2913,p2914,p2915,p2916,p2917,p2918,p2919,p2920,p2921,p2922,p2923,p2924,p2925,p2926,p2927,p2928,p2929,p2930,p2931,p2932,p2933,p2934,p2935,p2936,p2937,p2938,p2939,p2940,p2941,p2942,p2943,p2944,p2945,p2946,p2947,p2948,p2949,p2950,p2951,p2952,p2953,p2954,p2955,p2956,p2957,p2958,p2959,p2960,p2961,p2962,p2963,p2964,p2965,p2966,p2967,p2968,p2969,p2970,p2971,p2972,p2973,p2974,p2975,p2976,p2977,p2978,p2979,p2980,p2981,p2982,p2983,p2984,p2985,p2986,p2987,p2988,p2989,p2990,p2991,p2992,p2993,p2994,p2995,p2996,p2997,p2998,p2999,p3000,p3001,p3002,p3003,p3004,p3005,p3006,p3007,p3008,p3009,p3010,p3011,p3012,p3013,p3014,p3015,p3016,p3017,p3018,p3019,p3020,p3021,p3022,p3023,p3024,p3025,p3026,p3027,p3028,p3029,p3030,p3031,p3032,p3033,p3034,p3035,p3036,p3037,p3038,p3039,p3040,p3041,p3042,p3043,p3044,p3045,p3046,p3047,p3048,p3049,p3050,p3051,p3052,p3053,p3054,p3055,p3056,p3057,p3058,p3059,p3060,p3061,p3062,p3063,p3064,p3065,p3066,p3067,p3068,p3069,p3070,p3071,p3072,p3073,p3074,p3075,p3076,p3077,p3078,p3079,p3080,p3081,p3082,p3083,p3084,p3085,p3086,p3087,p3088,p3089,p3090,p3091,p3092,p3093,p3094,p3095,p3096,p3097,p3098,p3099,p3100,p3101,p3102,p3103,p3104,p3105,p3106,p3107,p3108,p3109,p3110,p3111,p3112,p3113,p3114,p3115,p3116,p3117,p3118,p3119,p3120,p3121,p3122,p3123,p3124,p3125,p3126,p3127,p3128,p3129,p3130,p3131,p3132,p3133,p3134,p3135,p3136,p3137,p3138,p3139,p3140,p3141,p3142,p3143,p3144,p3145,p3146,p3147,p3148,p3149,p3150,p3151,p3152,p3153,p3154,p3155,p3156,p3157,p3158,p3159,p3160,p3161,p3162,p3163,p3164,p3165,p3166,p3167,p3168,p3169,p3170,p3171,p3172,p3173,p3174,p3175,p3176,p3177,p3178,p3179,p3180,p3181,p3182,p3183,p3184,p3185,p3186,p3187,p3188,p3189,p3190,p3191,p3192,p3193,p3194,p3195,p3196,p3197,p3198,p3199,p3200,p3201,p3202,p3203,p3204,p3205,p3206,p3207,p3208,p3209,p3210,p3211,p3212,p3213,p3214,p3215,p3216,p3217,p3218,p3219,p3220,p3221,p3222,p3223,p3224,p3225,p3226,p3227,p3228,p3229,p3230,p3231,p3232,p3233,p3234,p3235,p3236,p3237,p3238,p3239,p3240,p3241,p3242,p3243,p3244,p3245,p3246,p3247,p3248,p3249,p3250,p3251,p3252,p3253,p3254,p3255,p3256,p3257,p3258,p3259,p3260,p3261,p3262,p3263,p3264,p3265,p3266,p3267,p3268,p3269,p3270,p3271,p3272,p3273,p3274,p3275,p3276,p3277,p3278,p3279,p3280,p3281,p3282,p3283,p3284,p3285,p3286,p3287,p3288,p3289,p3290,p3291,p3292,p3293,p3294,p3295,p3296,p3297,p3298,p3299,p3300,p3301,p3302,p3303,p3304,p3305,p3306,p3307,p3308,p3309,p3310,p3311,p3312,p3313,p3314,p3315,p3316,p3317,p3318,p3319,p3320,p3321,p3322,p3323,p3324,p3325,p3326,p3327,p3328,p3329,p3330,p3331,p3332,p3333,p3334,p3335,p3336,p3337,p3338,p3339,p3340,p3341,p3342,p3343,p3344,p3345,p3346,p3347,p3348,p3349,p3350,p3351,p3352,p3353,p3354,p3355,p3356,p3357,p3358,p3359,p3360,p3361,p3362,p3363,p3364,p3365,p3366,p3367,p3368,p3369,p3370,p3371,p3372,p3373,p3374,p3375,p3376,p3377,p3378,p3379,p3380,p3381,p3382,p3383,p3384,p3385,p3386,p3387,p3388,p3389,p3390,p3391,p3392,p3393,p3394,p3395,p3396,p3397,p3398,p3399,p3400,p3401,p3402,p3403,p3404,p3405,p3406,p3407,p3408,p3409,p3410,p3411,p3412,p3413,p3414,p3415,p3416,p3417,p3418,p3419,p3420,p3421,p3422,p3423,p3424,p3425,p3426,p3427,p3428,p3429,p3430,p3431,p3432,p3433,p3434,p3435,p3436,p3437,p3438,p3439,p3440,p3441,p3442,p3443,p3444,p3445,p3446,p3447,p3448,p3449,p3450,p3451,p3452,p3453,p3454,p3455,p3456,p3457,p3458,p3459,p3460,p3461,p3462,p3463,p3464,p3465,p3466,p3467,p3468,p3469,p3470,p3471,p3472,p3473,p3474,p3475,p3476,p3477,p3478,p3479,p3480,p3481,p3482,p3483,p3484,p3485,p3486,p3487,p3488,p3489,p3490,p3491,p3492,p3493,p3494,p3495,p3496,p3497,p3498,p3499,p3500,p3501,p3502,p3503,p3504,p3505,p3506,p3507,p3508,p3509,p3510,p3511,p3512,p3513,p3514,p3515,p3516,p3517,p3518,p3519,p3520,p3521,p3522,p3523,p3524,p3525,p3526,p3527,p3528,p3529,p3530,p3531,p3532,p3533,p3534,p3535,p3536,p3537,p3538,p3539,p3540,p3541,p3542,p3543,p3544,p3545,p3546,p3547,p3548,p3549,p3550,p3551,p3552,p3553,p3554,p3555,p3556,p3557,p3558,p3559,p3560,p3561,p3562,p3563,p3564,p3565,p3566,p3567,p3568,p3569,p3570,p3571,p3572,p3573,p3574,p3575,p3576,p3577,p3578,p3579,p3580,p3581,p3582,p3583,p3584,p3585,p3586,p3587,p3588,p3589,p3590,p3591,p3592,p3593,p3594,p3595,p3596,p3597,p3598,p3599,p3600,p3601,p3602,p3603,p3604,p3605,p3606,p3607,p3608,p3609,p3610,p3611,p3612,p3613,p3614,p3615,p3616,p3617,p3618,p3619,p3620,p3621,p3622,p3623,p3624,p3625,p3626,p3627,p3628,p3629,p3630,p3631,p3632,p3633,p3634,p3635,p3636,p3637,p3638,p3639,p3640,p3641,p3642,p3643,p3644,p3645,p3646,p3647,p3648,p3649,p3650,p3651,p3652,p3653,p3654,p3655,p3656,p3657,p3658,p3659,p3660,p3661,p3662,p3663,p3664,p3665,p3666,p3667,p3668,p3669,p3670,p3671,p3672,p3673,p3674,p3675,p3676,p3677,p3678,p3679,p3680,p3681,p3682,p3683,p3684,p3685,p3686,p3687,p3688,p3689,p3690,p3691,p3692,p3693,p3694,p3695,p3696,p3697,p3698,p3699,p3700,p3701,p3702,p3703,p3704,p3705,p3706,p3707,p3708,p3709,p3710,p3711,p3712,p3713,p3714,p3715,p3716,p3717,p3718,p3719,p3720,p3721,p3722,p3723,p3724,p3725,p3726,p3727,p3728,p3729,p3730,p3731,p3732,p3733,p3734,p3735,p3736,p3737,p3738,p3739,p3740,p3741,p3742,p3743,p3744,p3745,p3746,p3747,p3748,p3749,p3750,p3751,p3752,p3753,p3754,p3755,p3756,p3757,p3758,p3759,p3760,p3761,p3762,p3763,p3764,p3765,p3766,p3767,p3768,p3769,p3770,p3771,p3772,p3773,p3774,p3775,p3776,p3777,p3778,p3779,p3780,p3781,p3782,p3783,p3784,p3785,p3786,p3787,p3788,p3789,p3790,p3791,p3792,p3793,p3794,p3795,p3796,p3797,p3798,p3799,p3800,p3801,p3802,p3803,p3804,p3805,p3806,p3807,p3808,p3809,p3810,p3811,p3812,p3813,p3814,p3815,p3816,p3817,p3818,p3819,p3820,p3821,p3822,p3823,p3824,p3825,p3826,p3827,p3828,p3829,p3830,p3831,p3832,p3833,p3834,p3835,p3836,p3837,p3838,p3839,p3840,p3841,p3842,p3843,p3844,p3845,p3846,p3847,p3848,p3849,p3850,p3851,p3852,p3853,p3854,p3855,p3856,p3857,p3858,p3859,p3860,p3861,p3862,p3863,p3864,p3865,p3866,p3867,p3868,p3869,p3870,p3871,p3872,p3873,p3874,p3875,p3876,p3877,p3878,p3879,p3880,p3881,p3882,p3883,p3884,p3885,p3886,p3887,p3888,p3889,p3890,p3891,p3892,p3893,p3894,p3895,p3896,p3897,p3898,p3899,p3900,p3901,p3902,p3903,p3904,p3905,p3906,p3907,p3908,p3909,p3910,p3911,p3912,p3913,p3914,p3915,p3916,p3917,p3918,p3919,p3920,p3921,p3922,p3923,p3924,p3925,p3926,p3927,p3928,p3929,p3930,p3931,p3932,p3933,p3934,p3935,p3936,p3937,p3938,p3939,p3940,p3941,p3942,p3943,p3944,p3945,p3946,p3947,p3948,p3949,p3950,p3951,p3952,p3953,p3954,p3955,p3956,p3957,p3958,p3959,p3960,p3961,p3962,p3963,p3964,p3965,p3966,p3967,p3968,p3969,p3970,p3971,p3972,p3973,p3974,p3975,p3976,p3977,p3978,p3979,p3980,p3981,p3982,p3983,p3984,p3985,p3986,p3987,p3988,p3989,p3990,p3991,p3992,p3993,p3994,p3995,p3996,p3997,p3998,p3999,p4000,p4001,p4002,p4003,p4004,p4005,p4006,p4007,p4008,p4009,p4010,p4011,p4012,p4013,p4014,p4015,p4016,p4017,p4018,p4019,p4020,p4021,p4022,p4023,p4024,p4025,p4026,p4027,p4028,p4029,p4030,p4031,p4032,p4033,p4034,p4035,p4036,p4037,p4038,p4039,p4040,p4041,p4042,p4043,p4044,p4045,p4046,p4047,p4048,p4049,p4050,p4051,p4052,p4053,p4054,p4055,p4056,p4057,p4058,p4059,p4060,p4061,p4062,p4063,p4064,p4065,p4066,p4067,p4068,p4069,p4070,p4071,p4072,p4073,p4074,p4075,p4076,p4077,p4078,p4079,p4080,p4081,p4082,p4083,p4084,p4085,p4086,p4087,p4088,p4089,p4090,p4091,p4092,p4093,p4094,p4095,p4096,p4097,p4098,p4099,p4100,p4101,p4102,p4103,p4104,p4105,p4106,p4107,p4108,p4109,p4110,p4111,p4112,p4113,p4114,p4115,p4116,p4117,p4118,p4119,p4120,p4121,p4122,p4123,p4124,p4125,p4126,p4127,p4128,p4129,p4130,p4131,p4132,p4133,p4134,p4135,p4136,p4137,p4138,p4139,p4140,p4141,p4142,p4143,p4144,p4145,p4146,p4147,p4148,p4149,p4150,p4151,p4152,p4153,p4154,p4155,p4156,p4157,p4158,p4159,p4160,p4161,p4162,p4163,p4164,p4165,p4166,p4167,p4168,p4169,p4170,p4171,p4172,p4173,p4174,p4175,p4176,p4177,p4178,p4179,p4180,p4181,p4182,p4183,p4184,p4185,p4186,p4187,p4188,p4189,p4190,p4191,p4192,p4193,p4194,p4195,p4196,p4197,p4198,p4199,p4200,p4201,p4202,p4203,p4204,p4205,p4206,p4207,p4208,p4209,p4210,p4211,p4212,p4213,p4214,p4215,p4216,p4217,p4218,p4219,p4220,p4221,p4222,p4223,p4224,p4225,p4226,p4227,p4228,p4229,p4230,p4231,p4232,p4233,p4234,p4235,p4236,p4237,p4238,p4239,p4240,p4241,p4242,p4243,p4244,p4245,p4246,p4247,p4248,p4249,p4250,p4251,p4252,p4253,p4254,p4255,p4256,p4257,p4258,p4259,p4260,p4261,p4262,p4263,p4264,p4265,p4266,p4267,p4268,p4269,p4270,p4271,p4272,p4273,p4274,p4275,p4276,p4277,p4278,p4279,p4280,p4281,p4282,p4283,p4284,p4285,p4286,p4287,p4288,p4289,p4290,p4291,p4292,p4293,p4294,p4295,p4296,p4297,p4298,p4299,p4300,p4301,p4302,p4303,p4304,p4305,p4306,p4307,p4308,p4309,p4310,p4311,p4312,p4313,p4314,p4315,p4316,p4317,p4318,p4319,p4320,p4321,p4322,p4323,p4324,p4325,p4326,p4327,p4328,p4329,p4330,p4331,p4332,p4333,p4334,p4335,p4336,p4337,p4338,p4339,p4340,p4341,p4342,p4343,p4344,p4345,p4346,p4347,p4348,p4349,p4350,p4351,p4352,p4353,p4354,p4355,p4356,p4357,p4358,p4359,p4360,p4361,p4362,p4363,p4364,p4365,p4366,p4367,p4368,p4369,p4370,p4371,p4372,p4373,p4374,p4375,p4376,p4377,p4378,p4379,p4380,p4381,p4382,p4383,p4384,p4385,p4386,p4387,p4388,p4389,p4390,p4391,p4392,p4393,p4394,p4395,p4396,p4397,p4398,p4399,p4400,p4401,p4402,p4403,p4404,p4405,p4406,p4407,p4408,p4409,p4410,p4411,p4412,p4413,p4414,p4415,p4416,p4417,p4418,p4419,p4420,p4421,p4422,p4423,p4424,p4425,p4426,p4427,p4428,p4429,p4430,p4431,p4432,p4433,p4434,p4435,p4436,p4437,p4438,p4439,p4440,p4441,p4442,p4443,p4444,p4445,p4446,p4447,p4448,p4449,p4450,p4451,p4452,p4453,p4454,p4455,p4456,p4457,p4458,p4459,p4460,p4461,p4462,p4463,p4464,p4465,p4466,p4467,p4468,p4469,p4470,p4471,p4472,p4473,p4474,p4475,p4476,p4477,p4478,p4479,p4480,p4481,p4482,p4483,p4484,p4485,p4486,p4487,p4488,p4489,p4490,p4491,p4492,p4493,p4494,p4495,p4496,p4497,p4498,p4499,p4500,p4501,p4502,p4503,p4504,p4505,p4506,p4507,p4508,p4509,p4510,p4511,p4512,p4513,p4514,p4515,p4516,p4517,p4518,p4519,p4520,p4521,p4522,p4523,p4524,p4525,p4526,p4527,p4528,p4529,p4530,p4531,p4532,p4533,p4534,p4535,p4536,p4537,p4538,p4539,p4540,p4541,p4542,p4543,p4544,p4545,p4546,p4547,p4548,p4549,p4550,p4551,p4552,p4553,p4554,p4555,p4556,p4557,p4558,p4559,p4560,p4561,p4562,p4563,p4564,p4565,p4566,p4567,p4568,p4569,p4570,p4571,p4572,p4573,p4574,p4575,p4576,p4577,p4578,p4579,p4580,p4581,p4582,p4583,p4584,p4585,p4586,p4587,p4588,p4589,p4590,p4591,p4592,p4593,p4594,p4595,p4596,p4597,p4598,p4599,p4600,p4601,p4602,p4603,p4604,p4605,p4606,p4607,p4608,p4609,p4610,p4611,p4612,p4613,p4614,p4615,p4616,p4617,p4618,p4619,p4620,p4621,p4622,p4623,p4624,p4625,p4626,p4627,p4628,p4629,p4630,p4631,p4632,p4633,p4634,p4635,p4636,p4637,p4638,p4639,p4640,p4641,p4642,p4643,p4644,p4645,p4646,p4647,p4648,p4649,p4650,p4651,p4652,p4653,p4654,p4655,p4656,p4657,p4658,p4659,p4660,p4661,p4662,p4663,p4664,p4665,p4666,p4667,p4668,p4669,p4670,p4671,p4672,p4673,p4674,p4675,p4676,p4677,p4678,p4679,p4680,p4681,p4682,p4683,p4684,p4685,p4686,p4687,p4688,p4689,p4690,p4691,p4692,p4693,p4694,p4695,p4696,p4697,p4698,p4699,p4700,p4701,p4702,p4703,p4704,p4705,p4706,p4707,p4708,p4709,p4710,p4711,p4712,p4713,p4714,p4715,p4716,p4717,p4718,p4719,p4720,p4721,p4722,p4723,p4724,p4725,p4726,p4727,p4728,p4729,p4730,p4731,p4732,p4733,p4734,p4735,p4736,p4737,p4738,p4739,p4740,p4741,p4742,p4743,p4744,p4745,p4746,p4747,p4748,p4749,p4750,p4751,p4752,p4753,p4754,p4755,p4756,p4757,p4758,p4759,p4760,p4761,p4762,p4763,p4764,p4765,p4766,p4767,p4768,p4769,p4770,p4771,p4772,p4773,p4774,p4775,p4776,p4777,p4778,p4779,p4780,p4781,p4782,p4783,p4784,p4785,p4786,p4787,p4788,p4789,p4790,p4791,p4792,p4793,p4794,p4795,p4796,p4797,p4798,p4799,p4800,p4801,p4802,p4803,p4804,p4805,p4806,p4807,p4808,p4809,p4810,p4811,p4812,p4813,p4814,p4815,p4816,p4817,p4818,p4819,p4820,p4821,p4822,p4823,p4824,p4825,p4826,p4827,p4828,p4829,p4830,p4831,p4832,p4833,p4834,p4835,p4836,p4837,p4838,p4839,p4840,p4841,p4842,p4843,p4844,p4845,p4846,p4847,p4848,p4849,p4850,p4851,p4852,p4853,p4854,p4855,p4856,p4857,p4858,p4859,p4860,p4861,p4862,p4863,p4864,p4865,p4866,p4867,p4868,p4869,p4870,p4871,p4872,p4873,p4874,p4875,p4876,p4877,p4878,p4879,p4880,p4881,p4882,p4883,p4884,p4885,p4886,p4887,p4888,p4889,p4890,p4891,p4892,p4893,p4894,p4895,p4896,p4897,p4898,p4899,p4900,p4901,p4902,p4903,p4904,p4905,p4906,p4907,p4908,p4909,p4910,p4911,p4912,p4913,p4914,p4915,p4916,p4917,p4918,p4919,p4920,p4921,p4922,p4923,p4924,p4925,p4926,p4927,p4928,p4929,p4930,p4931,p4932,p4933,p4934,p4935,p4936,p4937,p4938,p4939,p4940,p4941,p4942,p4943,p4944,p4945,p4946,p4947,p4948,p4949,p4950,p4951,p4952,p4953,p4954,p4955,p4956,p4957,p4958,p4959,p4960,p4961,p4962,p4963,p4964,p4965,p4966,p4967,p4968,p4969,p4970,p4971,p4972,p4973,p4974,p4975,p4976,p4977,p4978,p4979,p4980,p4981,p4982,p4983,p4984,p4985,p4986,p4987,p4988,p4989,p4990,p4991,p4992,p4993,p4994,p4995,p4996,p4997,p4998,p4999,p5000,p5001,p5002,p5003,p5004,p5005,p5006,p5007,p5008,p5009,p5010,p5011,p5012,p5013,p5014,p5015,p5016,p5017,p5018,p5019,p5020,p5021,p5022,p5023,p5024,p5025,p5026,p5027,p5028,p5029,p5030,p5031,p5032,p5033,p5034,p5035,p5036,p5037,p5038,p5039,p5040,p5041,p5042,p5043,p5044,p5045,p5046,p5047,p5048,p5049,p5050,p5051,p5052,p5053,p5054,p5055,p5056,p5057,p5058,p5059,p5060,p5061,p5062,p5063,p5064,p5065,p5066,p5067,p5068,p5069,p5070,p5071,p5072,p5073,p5074,p5075,p5076,p5077,p5078,p5079,p5080,p5081,p5082,p5083,p5084,p5085,p5086,p5087,p5088,p5089,p5090,p5091,p5092,p5093,p5094,p5095,p5096,p5097,p5098,p5099,p5100,p5101,p5102,p5103,p5104,p5105,p5106,p5107,p5108,p5109,p5110,p5111,p5112,p5113,p5114,p5115,p5116,p5117,p5118,p5119,p5120,p5121,p5122,p5123,p5124,p5125,p5126,p5127,p5128,p5129,p5130,p5131,p5132,p5133,p5134,p5135,p5136,p5137,p5138,p5139,p5140,p5141,p5142,p5143,p5144,p5145,p5146,p5147,p5148,p5149,p5150,p5151,p5152,p5153,p5154,p5155,p5156,p5157,p5158,p5159,p5160,p5161,p5162,p5163,p5164,p5165,p5166,p5167,p5168,p5169,p5170,p5171,p5172,p5173,p5174,p5175,p5176,p5177,p5178,p5179,p5180,p5181,p5182,p5183,p5184,p5185,p5186,p5187,p5188,p5189,p5190,p5191,p5192,p5193,p5194,p5195,p5196,p5197,p5198,p5199,p5200,p5201,p5202,p5203,p5204,p5205,p5206,p5207,p5208,p5209,p5210,p5211,p5212,p5213,p5214,p5215,p5216,p5217,p5218,p5219,p5220,p5221,p5222,p5223,p5224,p5225,p5226,p5227,p5228,p5229,p5230,p5231,p5232,p5233,p5234,p5235,p5236,p5237,p5238,p5239,p5240,p5241,p5242,p5243,p5244,p5245,p5246,p5247,p5248,p5249,p5250,p5251,p5252,p5253,p5254,p5255,p5256,p5257,p5258,p5259,p5260,p5261,p5262,p5263,p5264,p5265,p5266,p5267,p5268,p5269,p5270,p5271,p5272,p5273,p5274,p5275,p5276,p5277,p5278,p5279,p5280,p5281,p5282,p5283,p5284,p5285,p5286,p5287,p5288,p5289,p5290,p5291,p5292,p5293,p5294,p5295,p5296,p5297,p5298,p5299,p5300,p5301,p5302,p5303,p5304,p5305,p5306,p5307,p5308,p5309,p5310,p5311,p5312,p5313,p5314,p5315,p5316,p5317,p5318,p5319,p5320,p5321,p5322,p5323,p5324,p5325,p5326,p5327,p5328,p5329,p5330,p5331,p5332,p5333,p5334,p5335,p5336,p5337,p5338,p5339,p5340,p5341,p5342,p5343,p5344,p5345,p5346,p5347,p5348,p5349,p5350,p5351,p5352,p5353,p5354,p5355,p5356,p5357,p5358,p5359,p5360,p5361,p5362,p5363,p5364,p5365,p5366,p5367,p5368,p5369,p5370,p5371,p5372,p5373,p5374,p5375,p5376,p5377,p5378,p5379,p5380,p5381,p5382,p5383,p5384,p5385,p5386,p5387,p5388,p5389,p5390,p5391,p5392,p5393,p5394,p5395,p5396,p5397,p5398,p5399,p5400,p5401,p5402,p5403,p5404,p5405,p5406,p5407,p5408,p5409,p5410,p5411,p5412,p5413,p5414,p5415,p5416,p5417,p5418,p5419,p5420,p5421,p5422,p5423,p5424,p5425,p5426,p5427,p5428,p5429,p5430,p5431,p5432,p5433,p5434,p5435,p5436,p5437,p5438,p5439,p5440,p5441,p5442,p5443,p5444,p5445,p5446,p5447,p5448,p5449,p5450,p5451,p5452,p5453,p5454,p5455,p5456,p5457,p5458,p5459,p5460,p5461,p5462,p5463,p5464,p5465,p5466,p5467,p5468,p5469,p5470,p5471,p5472,p5473,p5474,p5475,p5476,p5477,p5478,p5479,p5480,p5481,p5482,p5483,p5484,p5485,p5486,p5487,p5488,p5489,p5490,p5491,p5492,p5493,p5494,p5495,p5496,p5497,p5498,p5499,p5500,p5501,p5502,p5503,p5504,p5505,p5506,p5507,p5508,p5509,p5510,p5511,p5512,p5513,p5514,p5515,p5516,p5517,p5518,p5519,p5520,p5521,p5522,p5523,p5524,p5525,p5526,p5527,p5528,p5529,p5530,p5531,p5532,p5533,p5534,p5535,p5536,p5537,p5538,p5539,p5540,p5541,p5542,p5543,p5544,p5545,p5546,p5547,p5548,p5549,p5550,p5551,p5552,p5553,p5554,p5555,p5556,p5557,p5558,p5559,p5560,p5561,p5562,p5563,p5564,p5565,p5566,p5567,p5568,p5569,p5570,p5571,p5572,p5573,p5574,p5575,p5576,p5577,p5578,p5579,p5580,p5581,p5582,p5583,p5584,p5585,p5586,p5587,p5588,p5589,p5590,p5591,p5592,p5593,p5594,p5595,p5596,p5597,p5598,p5599,p5600,p5601,p5602,p5603,p5604,p5605,p5606,p5607,p5608,p5609,p5610,p5611,p5612,p5613,p5614,p5615,p5616,p5617,p5618,p5619,p5620,p5621,p5622,p5623,p5624,p5625,p5626,p5627,p5628,p5629,p5630,p5631,p5632,p5633,p5634,p5635,p5636,p5637,p5638,p5639,p5640,p5641,p5642,p5643,p5644,p5645,p5646,p5647,p5648,p5649,p5650,p5651,p5652,p5653,p5654,p5655,p5656,p5657,p5658,p5659,p5660,p5661,p5662,p5663,p5664,p5665,p5666,p5667,p5668,p5669,p5670,p5671,p5672,p5673,p5674,p5675,p5676,p5677,p5678,p5679,p5680,p5681,p5682,p5683,p5684,p5685,p5686,p5687,p5688,p5689,p5690,p5691,p5692,p5693,p5694,p5695,p5696,p5697,p5698,p5699,p5700,p5701,p5702,p5703,p5704,p5705,p5706,p5707,p5708,p5709,p5710,p5711,p5712,p5713,p5714,p5715,p5716,p5717,p5718,p5719,p5720,p5721,p5722,p5723,p5724,p5725,p5726,p5727,p5728,p5729,p5730,p5731,p5732,p5733,p5734,p5735,p5736,p5737,p5738,p5739,p5740,p5741,p5742,p5743,p5744,p5745,p5746,p5747,p5748,p5749,p5750,p5751,p5752,p5753,p5754,p5755,p5756,p5757,p5758,p5759,p5760,p5761,p5762,p5763,p5764,p5765,p5766,p5767,p5768,p5769,p5770,p5771,p5772,p5773,p5774,p5775,p5776,p5777,p5778,p5779,p5780,p5781,p5782,p5783,p5784,p5785,p5786,p5787,p5788,p5789,p5790,p5791,p5792,p5793,p5794,p5795,p5796,p5797,p5798,p5799,p5800,p5801,p5802,p5803,p5804,p5805,p5806,p5807,p5808,p5809,p5810,p5811,p5812,p5813,p5814,p5815,p5816,p5817,p5818,p5819,p5820,p5821,p5822,p5823,p5824,p5825,p5826,p5827,p5828,p5829,p5830,p5831,p5832,p5833,p5834,p5835,p5836,p5837,p5838,p5839,p5840,p5841,p5842,p5843,p5844,p5845,p5846,p5847,p5848,p5849,p5850,p5851,p5852,p5853,p5854,p5855,p5856,p5857,p5858,p5859,p5860,p5861,p5862,p5863,p5864,p5865,p5866,p5867,p5868,p5869,p5870,p5871,p5872,p5873,p5874,p5875,p5876,p5877,p5878,p5879,p5880,p5881,p5882,p5883,p5884,p5885,p5886,p5887,p5888,p5889,p5890,p5891,p5892,p5893,p5894,p5895,p5896,p5897,p5898,p5899,p5900,p5901,p5902,p5903,p5904,p5905,p5906,p5907,p5908,p5909,p5910,p5911,p5912,p5913,p5914,p5915,p5916,p5917,p5918,p5919,p5920,p5921,p5922,p5923,p5924,p5925,p5926,p5927,p5928,p5929,p5930,p5931,p5932,p5933,p5934,p5935,p5936,p5937,p5938,p5939,p5940,p5941,p5942,p5943,p5944,p5945,p5946,p5947,p5948,p5949,p5950,p5951,p5952,p5953,p5954,p5955,p5956,p5957,p5958,p5959,p5960,p5961,p5962,p5963,p5964,p5965,p5966,p5967,p5968,p5969,p5970,p5971,p5972,p5973,p5974,p5975,p5976,p5977,p5978,p5979,p5980,p5981,p5982,p5983,p5984,p5985,p5986,p5987,p5988,p5989,p5990,p5991,p5992,p5993,p5994,p5995,p5996,p5997,p5998,p5999,p6000,p6001,p6002,p6003,p6004,p6005,p6006,p6007,p6008,p6009,p6010,p6011,p6012,p6013,p6014,p6015,p6016,p6017,p6018,p6019,p6020,p6021,p6022,p6023,p6024,p6025,p6026,p6027,p6028,p6029,p6030,p6031,p6032,p6033,p6034,p6035,p6036,p6037,p6038,p6039,p6040,p6041,p6042,p6043,p6044,p6045,p6046,p6047,p6048,p6049,p6050,p6051,p6052,p6053,p6054,p6055,p6056,p6057,p6058,p6059,p6060,p6061,p6062,p6063,p6064,p6065,p6066,p6067,p6068,p6069,p6070,p6071,p6072,p6073,p6074,p6075,p6076,p6077,p6078,p6079,p6080,p6081,p6082,p6083,p6084,p6085,p6086,p6087,p6088,p6089,p6090,p6091,p6092,p6093,p6094,p6095,p6096,p6097,p6098,p6099,p6100,p6101,p6102,p6103,p6104,p6105,p6106,p6107,p6108,p6109,p6110,p6111,p6112,p6113,p6114,p6115,p6116,p6117,p6118,p6119,p6120,p6121,p6122,p6123,p6124,p6125,p6126,p6127,p6128,p6129,p6130,p6131,p6132,p6133,p6134,p6135,p6136,p6137,p6138,p6139,p6140,p6141,p6142,p6143,p6144,p6145,p6146,p6147,p6148,p6149,p6150,p6151,p6152,p6153,p6154,p6155,p6156,p6157,p6158,p6159,p6160,p6161,p6162,p6163,p6164,p6165,p6166,p6167,p6168,p6169,p6170,p6171,p6172,p6173,p6174,p6175,p6176,p6177,p6178,p6179,p6180,p6181,p6182,p6183,p6184,p6185,p6186,p6187,p6188,p6189,p6190,p6191,p6192,p6193,p6194,p6195,p6196,p6197,p6198,p6199,p6200,p6201,p6202,p6203,p6204,p6205,p6206,p6207,p6208,p6209,p6210,p6211,p6212,p6213,p6214,p6215,p6216,p6217,p6218,p6219,p6220,p6221,p6222,p6223,p6224,p6225,p6226,p6227,p6228,p6229,p6230,p6231,p6232,p6233,p6234,p6235,p6236,p6237,p6238,p6239,p6240,p6241,p6242,p6243,p6244,p6245,p6246,p6247,p6248,p6249,p6250,p6251,p6252,p6253,p6254,p6255,p6256,p6257,p6258,p6259,p6260,p6261,p6262,p6263,p6264,p6265,p6266,p6267,p6268,p6269,p6270,p6271,p6272,p6273,p6274,p6275,p6276,p6277,p6278,p6279,p6280,p6281,p6282,p6283,p6284,p6285,p6286,p6287,p6288,p6289,p6290,p6291,p6292,p6293,p6294,p6295,p6296,p6297,p6298,p6299,p6300,p6301,p6302,p6303,p6304,p6305,p6306,p6307,p6308,p6309,p6310,p6311,p6312,p6313,p6314,p6315,p6316,p6317,p6318,p6319,p6320,p6321,p6322,p6323,p6324,p6325,p6326,p6327,p6328,p6329,p6330,p6331,p6332,p6333,p6334,p6335,p6336,p6337,p6338,p6339,p6340,p6341,p6342,p6343,p6344,p6345,p6346,p6347,p6348,p6349,p6350,p6351,p6352,p6353,p6354,p6355,p6356,p6357,p6358,p6359,p6360,p6361,p6362,p6363,p6364,p6365,p6366,p6367,p6368,p6369,p6370,p6371,p6372,p6373,p6374,p6375,p6376,p6377,p6378,p6379,p6380,p6381,p6382,p6383,p6384,p6385,p6386,p6387,p6388,p6389,p6390,p6391,p6392,p6393,p6394,p6395,p6396,p6397,p6398,p6399,p6400,p6401,p6402,p6403,p6404,p6405,p6406,p6407,p6408,p6409,p6410,p6411,p6412,p6413,p6414,p6415,p6416,p6417,p6418,p6419,p6420,p6421,p6422,p6423,p6424,p6425,p6426,p6427,p6428,p6429,p6430,p6431,p6432,p6433,p6434,p6435,p6436,p6437,p6438,p6439,p6440,p6441,p6442,p6443,p6444,p6445,p6446,p6447,p6448,p6449,p6450,p6451,p6452,p6453,p6454,p6455,p6456,p6457,p6458,p6459,p6460,p6461,p6462,p6463,p6464,p6465,p6466,p6467,p6468,p6469,p6470,p6471,p6472,p6473,p6474,p6475,p6476,p6477,p6478,p6479,p6480,p6481,p6482,p6483,p6484,p6485,p6486,p6487,p6488,p6489,p6490,p6491,p6492,p6493,p6494,p6495,p6496,p6497,p6498,p6499,p6500,p6501,p6502,p6503,p6504,p6505,p6506,p6507,p6508,p6509,p6510,p6511,p6512,p6513,p6514,p6515,p6516,p6517,p6518,p6519,p6520,p6521,p6522,p6523,p6524,p6525,p6526,p6527,p6528,p6529,p6530,p6531,p6532,p6533,p6534,p6535,p6536,p6537,p6538,p6539,p6540,p6541,p6542,p6543,p6544,p6545,p6546,p6547,p6548,p6549,p6550,p6551,p6552,p6553,p6554,p6555,p6556,p6557,p6558,p6559,p6560,p6561,p6562,p6563,p6564,p6565,p6566,p6567,p6568,p6569,p6570,p6571,p6572,p6573,p6574,p6575,p6576,p6577,p6578,p6579,p6580,p6581,p6582,p6583,p6584,p6585,p6586,p6587,p6588,p6589,p6590,p6591,p6592,p6593,p6594,p6595,p6596,p6597,p6598,p6599,p6600,p6601,p6602,p6603,p6604,p6605,p6606,p6607,p6608,p6609,p6610,p6611,p6612,p6613,p6614,p6615,p6616,p6617,p6618,p6619,p6620,p6621,p6622,p6623,p6624,p6625,p6626,p6627,p6628,p6629,p6630,p6631,p6632,p6633,p6634,p6635,p6636,p6637,p6638,p6639,p6640,p6641,p6642,p6643,p6644,p6645,p6646,p6647,p6648,p6649,p6650,p6651,p6652,p6653,p6654,p6655,p6656,p6657,p6658,p6659,p6660,p6661,p6662,p6663,p6664,p6665,p6666,p6667,p6668,p6669,p6670,p6671,p6672,p6673,p6674,p6675,p6676,p6677,p6678,p6679,p6680,p6681,p6682,p6683,p6684,p6685,p6686,p6687,p6688,p6689,p6690,p6691,p6692,p6693,p6694,p6695,p6696,p6697,p6698,p6699,p6700,p6701,p6702,p6703,p6704,p6705,p6706,p6707,p6708,p6709,p6710,p6711,p6712,p6713,p6714,p6715,p6716,p6717,p6718,p6719,p6720,p6721,p6722,p6723,p6724,p6725,p6726,p6727,p6728,p6729,p6730,p6731,p6732,p6733,p6734,p6735,p6736,p6737,p6738,p6739,p6740,p6741,p6742,p6743,p6744,p6745,p6746,p6747,p6748,p6749,p6750,p6751,p6752,p6753,p6754,p6755,p6756,p6757,p6758,p6759,p6760,p6761,p6762,p6763,p6764,p6765,p6766,p6767,p6768,p6769,p6770,p6771,p6772,p6773,p6774,p6775,p6776,p6777,p6778,p6779,p6780,p6781,p6782,p6783,p6784,p6785,p6786,p6787,p6788,p6789,p6790,p6791,p6792,p6793,p6794,p6795,p6796,p6797,p6798,p6799,p6800,p6801,p6802,p6803,p6804,p6805,p6806,p6807,p6808,p6809,p6810,p6811,p6812,p6813,p6814,p6815,p6816,p6817,p6818,p6819,p6820,p6821,p6822,p6823,p6824,p6825,p6826,p6827,p6828,p6829,p6830,p6831,p6832,p6833,p6834,p6835,p6836,p6837,p6838,p6839,p6840,p6841,p6842,p6843,p6844,p6845,p6846,p6847,p6848,p6849,p6850,p6851,p6852,p6853,p6854,p6855,p6856,p6857,p6858,p6859,p6860,p6861,p6862,p6863,p6864,p6865,p6866,p6867,p6868,p6869,p6870,p6871,p6872,p6873,p6874,p6875,p6876,p6877,p6878,p6879,p6880,p6881,p6882,p6883,p6884,p6885,p6886,p6887,p6888,p6889,p6890,p6891,p6892,p6893,p6894,p6895,p6896,p6897,p6898,p6899,p6900,p6901,p6902,p6903,p6904,p6905,p6906,p6907,p6908,p6909,p6910,p6911,p6912,p6913,p6914,p6915,p6916,p6917,p6918,p6919,p6920,p6921,p6922,p6923,p6924,p6925,p6926,p6927,p6928,p6929,p6930,p6931,p6932,p6933,p6934,p6935,p6936,p6937,p6938,p6939,p6940,p6941,p6942,p6943,p6944,p6945,p6946,p6947,p6948,p6949,p6950,p6951,p6952,p6953,p6954,p6955,p6956,p6957,p6958,p6959,p6960,p6961,p6962,p6963,p6964,p6965,p6966,p6967,p6968,p6969,p6970,p6971,p6972,p6973,p6974,p6975,p6976,p6977,p6978,p6979,p6980,p6981,p6982,p6983,p6984,p6985,p6986,p6987,p6988,p6989,p6990,p6991,p6992,p6993,p6994,p6995,p6996,p6997,p6998,p6999,p7000,p7001,p7002,p7003,p7004,p7005,p7006,p7007,p7008,p7009,p7010,p7011,p7012,p7013,p7014,p7015,p7016,p7017,p7018,p7019,p7020,p7021,p7022,p7023,p7024,p7025,p7026,p7027,p7028,p7029,p7030,p7031,p7032,p7033,p7034,p7035,p7036,p7037,p7038,p7039,p7040,p7041,p7042,p7043,p7044,p7045,p7046,p7047,p7048,p7049,p7050,p7051,p7052,p7053,p7054,p7055,p7056,p7057,p7058,p7059,p7060,p7061,p7062,p7063,p7064,p7065,p7066,p7067,p7068,p7069,p7070,p7071,p7072,p7073,p7074,p7075,p7076,p7077,p7078,p7079,p7080,p7081,p7082,p7083,p7084,p7085,p7086,p7087,p7088,p7089,p7090,p7091,p7092,p7093,p7094,p7095,p7096,p7097,p7098,p7099,p7100,p7101,p7102,p7103,p7104,p7105,p7106,p7107,p7108,p7109,p7110,p7111,p7112,p7113,p7114,p7115,p7116,p7117,p7118,p7119,p7120,p7121,p7122,p7123,p7124,p7125,p7126,p7127,p7128,p7129,p7130,p7131,p7132,p7133,p7134,p7135,p7136,p7137,p7138,p7139,p7140,p7141,p7142,p7143,p7144,p7145,p7146,p7147,p7148,p7149,p7150,p7151,p7152,p7153,p7154,p7155,p7156,p7157,p7158,p7159,p7160,p7161,p7162,p7163,p7164,p7165,p7166,p7167,p7168,p7169,p7170,p7171,p7172,p7173,p7174,p7175,p7176,p7177,p7178,p7179,p7180,p7181,p7182,p7183,p7184,p7185,p7186,p7187,p7188,p7189,p7190,p7191,p7192,p7193,p7194,p7195,p7196,p7197,p7198,p7199,p7200,p7201,p7202,p7203,p7204,p7205,p7206,p7207,p7208,p7209,p7210,p7211,p7212,p7213,p7214,p7215,p7216,p7217,p7218,p7219,p7220,p7221,p7222,p7223,p7224,p7225,p7226,p7227,p7228,p7229,p7230,p7231,p7232,p7233,p7234,p7235,p7236,p7237,p7238,p7239,p7240,p7241,p7242,p7243,p7244,p7245,p7246,p7247,p7248,p7249,p7250,p7251,p7252,p7253,p7254,p7255,p7256,p7257,p7258,p7259,p7260,p7261,p7262,p7263,p7264,p7265,p7266,p7267,p7268,p7269,p7270,p7271,p7272,p7273,p7274,p7275,p7276,p7277,p7278,p7279,p7280,p7281,p7282,p7283,p7284,p7285,p7286,p7287,p7288,p7289,p7290,p7291,p7292,p7293,p7294,p7295,p7296,p7297,p7298,p7299,p7300,p7301,p7302,p7303,p7304,p7305,p7306,p7307,p7308,p7309,p7310,p7311,p7312,p7313,p7314,p7315,p7316,p7317,p7318,p7319,p7320,p7321,p7322,p7323,p7324,p7325,p7326,p7327,p7328,p7329,p7330,p7331,p7332,p7333,p7334,p7335,p7336,p7337,p7338,p7339,p7340,p7341,p7342,p7343,p7344,p7345,p7346,p7347,p7348,p7349,p7350,p7351,p7352,p7353,p7354,p7355,p7356,p7357,p7358,p7359,p7360,p7361,p7362,p7363,p7364,p7365,p7366,p7367,p7368,p7369,p7370,p7371,p7372,p7373,p7374,p7375,p7376,p7377,p7378,p7379,p7380,p7381,p7382,p7383,p7384,p7385,p7386,p7387,p7388,p7389,p7390,p7391,p7392,p7393,p7394,p7395,p7396,p7397,p7398,p7399,p7400,p7401,p7402,p7403,p7404,p7405,p7406,p7407,p7408,p7409,p7410,p7411,p7412,p7413,p7414,p7415,p7416,p7417,p7418,p7419,p7420,p7421,p7422,p7423,p7424,p7425,p7426,p7427,p7428,p7429,p7430,p7431,p7432,p7433,p7434,p7435,p7436,p7437,p7438,p7439,p7440,p7441,p7442,p7443,p7444,p7445,p7446,p7447,p7448,p7449,p7450,p7451,p7452,p7453,p7454,p7455,p7456,p7457,p7458,p7459,p7460,p7461,p7462,p7463,p7464,p7465,p7466,p7467,p7468,p7469,p7470,p7471,p7472,p7473,p7474,p7475,p7476,p7477,p7478,p7479,p7480,p7481,p7482,p7483,p7484,p7485,p7486,p7487,p7488,p7489,p7490,p7491,p7492,p7493,p7494,p7495,p7496,p7497,p7498,p7499,p7500,p7501,p7502,p7503,p7504,p7505,p7506,p7507,p7508,p7509,p7510,p7511,p7512,p7513,p7514,p7515,p7516,p7517,p7518,p7519,p7520,p7521,p7522,p7523,p7524,p7525,p7526,p7527,p7528,p7529,p7530,p7531,p7532,p7533,p7534,p7535,p7536,p7537,p7538,p7539,p7540,p7541,p7542,p7543,p7544,p7545,p7546,p7547,p7548,p7549,p7550,p7551,p7552,p7553,p7554,p7555,p7556,p7557,p7558,p7559,p7560,p7561,p7562,p7563,p7564,p7565,p7566,p7567,p7568,p7569,p7570,p7571,p7572,p7573,p7574,p7575,p7576,p7577,p7578,p7579,p7580,p7581,p7582,p7583,p7584,p7585,p7586,p7587,p7588,p7589,p7590,p7591,p7592,p7593,p7594,p7595,p7596,p7597,p7598,p7599,p7600,p7601,p7602,p7603,p7604,p7605,p7606,p7607,p7608,p7609,p7610,p7611,p7612,p7613,p7614,p7615,p7616,p7617,p7618,p7619,p7620,p7621,p7622,p7623,p7624,p7625,p7626,p7627,p7628,p7629,p7630,p7631,p7632,p7633,p7634,p7635,p7636,p7637,p7638,p7639,p7640,p7641,p7642,p7643,p7644,p7645,p7646,p7647,p7648,p7649,p7650,p7651,p7652,p7653,p7654,p7655,p7656,p7657,p7658,p7659,p7660,p7661,p7662,p7663,p7664,p7665,p7666,p7667,p7668,p7669,p7670,p7671,p7672,p7673,p7674,p7675,p7676,p7677,p7678,p7679,p7680,p7681,p7682,p7683,p7684,p7685,p7686,p7687,p7688,p7689,p7690,p7691,p7692,p7693,p7694,p7695,p7696,p7697,p7698,p7699,p7700,p7701,p7702,p7703,p7704,p7705,p7706,p7707,p7708,p7709,p7710,p7711,p7712,p7713,p7714,p7715,p7716,p7717,p7718,p7719,p7720,p7721,p7722,p7723,p7724,p7725,p7726,p7727,p7728,p7729,p7730,p7731,p7732,p7733,p7734,p7735,p7736,p7737,p7738,p7739,p7740,p7741,p7742,p7743,p7744,p7745,p7746,p7747,p7748,p7749,p7750,p7751,p7752,p7753,p7754,p7755,p7756,p7757,p7758,p7759,p7760,p7761,p7762,p7763,p7764,p7765,p7766,p7767,p7768,p7769,p7770,p7771,p7772,p7773,p7774,p7775,p7776,p7777,p7778,p7779,p7780,p7781,p7782,p7783,p7784,p7785,p7786,p7787,p7788,p7789,p7790,p7791,p7792,p7793,p7794,p7795,p7796,p7797,p7798,p7799,p7800,p7801,p7802,p7803,p7804,p7805,p7806,p7807,p7808,p7809,p7810,p7811,p7812,p7813,p7814,p7815,p7816,p7817,p7818,p7819,p7820,p7821,p7822,p7823,p7824,p7825,p7826,p7827,p7828,p7829,p7830,p7831,p7832,p7833,p7834,p7835,p7836,p7837,p7838,p7839,p7840,p7841,p7842,p7843,p7844,p7845,p7846,p7847,p7848,p7849,p7850,p7851,p7852,p7853,p7854,p7855,p7856,p7857,p7858,p7859,p7860,p7861,p7862,p7863,p7864,p7865,p7866,p7867,p7868,p7869,p7870,p7871,p7872,p7873,p7874,p7875,p7876,p7877,p7878,p7879,p7880,p7881,p7882,p7883,p7884,p7885,p7886,p7887,p7888,p7889,p7890,p7891,p7892,p7893,p7894,p7895,p7896,p7897,p7898,p7899,p7900,p7901,p7902,p7903,p7904,p7905,p7906,p7907,p7908,p7909,p7910,p7911,p7912,p7913,p7914,p7915,p7916,p7917,p7918,p7919,p7920,p7921,p7922,p7923,p7924,p7925,p7926,p7927,p7928,p7929,p7930,p7931,p7932,p7933,p7934,p7935,p7936,p7937,p7938,p7939,p7940,p7941,p7942,p7943,p7944,p7945,p7946,p7947,p7948,p7949,p7950,p7951,p7952,p7953,p7954,p7955,p7956,p7957,p7958,p7959,p7960,p7961,p7962,p7963,p7964,p7965,p7966,p7967,p7968,p7969,p7970,p7971,p7972,p7973,p7974,p7975,p7976,p7977,p7978,p7979,p7980,p7981,p7982,p7983,p7984,p7985,p7986,p7987,p7988,p7989,p7990,p7991,p7992,p7993,p7994,p7995,p7996,p7997,p7998,p7999,p8000,p8001,p8002,p8003,p8004,p8005,p8006,p8007,p8008,p8009,p8010,p8011,p8012,p8013,p8014,p8015,p8016,p8017,p8018,p8019,p8020,p8021,p8022,p8023,p8024,p8025,p8026,p8027,p8028,p8029,p8030,p8031,p8032,p8033,p8034,p8035,p8036,p8037,p8038,p8039,p8040,p8041,p8042,p8043,p8044,p8045,p8046,p8047,p8048,p8049,p8050,p8051,p8052,p8053,p8054,p8055,p8056,p8057,p8058,p8059,p8060,p8061,p8062,p8063,p8064,p8065,p8066,p8067,p8068,p8069,p8070,p8071,p8072,p8073,p8074,p8075,p8076,p8077,p8078,p8079,p8080,p8081,p8082,p8083,p8084,p8085,p8086,p8087,p8088,p8089,p8090,p8091,p8092,p8093,p8094,p8095,p8096,p8097,p8098,p8099,p8100,p8101,p8102,p8103,p8104,p8105,p8106,p8107,p8108,p8109,p8110,p8111,p8112,p8113,p8114,p8115,p8116,p8117,p8118,p8119,p8120,p8121,p8122,p8123,p8124,p8125,p8126,p8127,p8128,p8129,p8130,p8131,p8132,p8133,p8134,p8135,p8136,p8137,p8138,p8139,p8140,p8141,p8142,p8143,p8144,p8145,p8146,p8147,p8148,p8149,p8150,p8151,p8152,p8153,p8154,p8155,p8156,p8157,p8158,p8159,p8160,p8161,p8162,p8163,p8164,p8165,p8166,p8167,p8168,p8169,p8170,p8171,p8172,p8173,p8174,p8175,p8176,p8177,p8178,p8179,p8180,p8181,p8182,p8183,p8184,p8185,p8186,p8187,p8188,p8189,p8190,p8191,p8192,p8193,p8194,p8195,p8196,p8197,p8198,p8199,p8200,p8201,p8202,p8203,p8204,p8205,p8206,p8207,p8208,p8209,p8210,p8211,p8212,p8213,p8214,p8215,p8216,p8217,p8218,p8219,p8220,p8221,p8222,p8223,p8224,p8225,p8226,p8227,p8228,p8229,p8230,p8231,p8232,p8233,p8234,p8235,p8236,p8237,p8238,p8239,p8240,p8241,p8242,p8243,p8244,p8245,p8246,p8247,p8248,p8249,p8250,p8251,p8252,p8253,p8254,p8255,p8256,p8257,p8258,p8259,p8260,p8261,p8262,p8263,p8264,p8265,p8266,p8267,p8268,p8269,p8270,p8271,p8272,p8273,p8274,p8275,p8276,p8277,p8278,p8279,p8280,p8281,p8282,p8283,p8284,p8285,p8286,p8287,p8288,p8289,p8290,p8291,p8292,p8293,p8294,p8295,p8296,p8297,p8298,p8299,p8300,p8301,p8302,p8303,p8304,p8305,p8306,p8307,p8308,p8309,p8310,p8311,p8312,p8313,p8314,p8315,p8316,p8317,p8318,p8319,p8320,p8321,p8322,p8323,p8324,p8325,p8326,p8327,p8328,p8329,p8330,p8331,p8332,p8333,p8334,p8335,p8336,p8337,p8338,p8339,p8340,p8341,p8342,p8343,p8344,p8345,p8346,p8347,p8348,p8349,p8350,p8351,p8352,p8353,p8354,p8355,p8356,p8357,p8358,p8359,p8360,p8361,p8362,p8363,p8364,p8365,p8366,p8367,p8368,p8369,p8370,p8371,p8372,p8373,p8374,p8375,p8376,p8377,p8378,p8379,p8380,p8381,p8382,p8383,p8384,p8385,p8386,p8387,p8388,p8389,p8390,p8391,p8392,p8393,p8394,p8395,p8396,p8397,p8398,p8399,p8400,p8401,p8402,p8403,p8404,p8405,p8406,p8407,p8408,p8409,p8410,p8411,p8412,p8413,p8414,p8415,p8416,p8417,p8418,p8419,p8420,p8421,p8422,p8423,p8424,p8425,p8426,p8427,p8428,p8429,p8430,p8431,p8432,p8433,p8434,p8435,p8436,p8437,p8438,p8439,p8440,p8441,p8442,p8443,p8444,p8445,p8446,p8447,p8448,p8449,p8450,p8451,p8452,p8453,p8454,p8455,p8456,p8457,p8458,p8459,p8460,p8461,p8462,p8463,p8464,p8465,p8466,p8467,p8468,p8469,p8470,p8471,p8472,p8473,p8474,p8475,p8476,p8477,p8478,p8479,p8480,p8481,p8482,p8483,p8484,p8485,p8486,p8487,p8488,p8489,p8490,p8491,p8492,p8493,p8494,p8495,p8496,p8497,p8498,p8499,p8500,p8501,p8502,p8503,p8504,p8505,p8506,p8507,p8508,p8509,p8510,p8511,p8512,p8513,p8514,p8515,p8516,p8517,p8518,p8519,p8520,p8521,p8522,p8523,p8524,p8525,p8526,p8527,p8528,p8529,p8530,p8531,p8532,p8533,p8534,p8535,p8536,p8537,p8538,p8539,p8540,p8541,p8542,p8543,p8544,p8545,p8546,p8547,p8548,p8549,p8550,p8551,p8552,p8553,p8554,p8555,p8556,p8557,p8558,p8559,p8560,p8561,p8562,p8563,p8564,p8565,p8566,p8567,p8568,p8569,p8570,p8571,p8572,p8573,p8574,p8575,p8576,p8577,p8578,p8579,p8580,p8581,p8582,p8583,p8584,p8585,p8586,p8587,p8588,p8589,p8590,p8591,p8592,p8593,p8594,p8595,p8596,p8597,p8598,p8599,p8600,p8601,p8602,p8603,p8604,p8605,p8606,p8607,p8608,p8609,p8610,p8611,p8612,p8613,p8614,p8615,p8616,p8617,p8618,p8619,p8620,p8621,p8622,p8623,p8624,p8625,p8626,p8627,p8628,p8629,p8630,p8631,p8632,p8633,p8634,p8635,p8636,p8637,p8638,p8639,p8640,p8641,p8642,p8643,p8644,p8645,p8646,p8647,p8648,p8649,p8650,p8651,p8652,p8653,p8654,p8655,p8656,p8657,p8658,p8659,p8660,p8661,p8662,p8663,p8664,p8665,p8666,p8667,p8668,p8669,p8670,p8671,p8672,p8673,p8674,p8675,p8676,p8677,p8678,p8679,p8680,p8681,p8682,p8683,p8684,p8685,p8686,p8687,p8688,p8689,p8690,p8691,p8692,p8693,p8694,p8695,p8696,p8697,p8698,p8699,p8700,p8701,p8702,p8703,p8704,p8705,p8706,p8707,p8708,p8709,p8710,p8711,p8712,p8713,p8714,p8715,p8716,p8717,p8718,p8719,p8720,p8721,p8722,p8723,p8724,p8725,p8726,p8727,p8728,p8729,p8730,p8731,p8732,p8733,p8734,p8735,p8736,p8737,p8738,p8739,p8740,p8741,p8742,p8743,p8744,p8745,p8746,p8747,p8748,p8749,p8750,p8751,p8752,p8753,p8754,p8755,p8756,p8757,p8758,p8759,p8760,p8761,p8762,p8763,p8764,p8765,p8766,p8767,p8768,p8769,p8770,p8771,p8772,p8773,p8774,p8775,p8776,p8777,p8778,p8779,p8780,p8781,p8782,p8783,p8784,p8785,p8786,p8787,p8788,p8789,p8790,p8791,p8792,p8793,p8794,p8795,p8796,p8797,p8798,p8799,p8800,p8801,p8802,p8803,p8804,p8805,p8806,p8807,p8808,p8809,p8810,p8811,p8812,p8813,p8814,p8815,p8816,p8817,p8818,p8819,p8820,p8821,p8822,p8823,p8824,p8825,p8826,p8827,p8828,p8829,p8830,p8831,p8832,p8833,p8834,p8835,p8836,p8837,p8838,p8839,p8840,p8841,p8842,p8843,p8844,p8845,p8846,p8847,p8848,p8849,p8850,p8851,p8852,p8853,p8854,p8855,p8856,p8857,p8858,p8859,p8860,p8861,p8862,p8863,p8864,p8865,p8866,p8867,p8868,p8869,p8870,p8871,p8872,p8873,p8874,p8875,p8876,p8877,p8878,p8879,p8880,p8881,p8882,p8883,p8884,p8885,p8886,p8887,p8888,p8889,p8890,p8891,p8892,p8893,p8894,p8895,p8896,p8897,p8898,p8899,p8900,p8901,p8902,p8903,p8904,p8905,p8906,p8907,p8908,p8909,p8910,p8911,p8912,p8913,p8914,p8915,p8916,p8917,p8918,p8919,p8920,p8921,p8922,p8923,p8924,p8925,p8926,p8927,p8928,p8929,p8930,p8931,p8932,p8933,p8934,p8935,p8936,p8937,p8938,p8939,p8940,p8941,p8942,p8943,p8944,p8945,p8946,p8947,p8948,p8949,p8950,p8951,p8952,p8953,p8954,p8955,p8956,p8957,p8958,p8959,p8960,p8961,p8962,p8963,p8964,p8965,p8966,p8967,p8968,p8969,p8970,p8971,p8972,p8973,p8974,p8975,p8976,p8977,p8978,p8979,p8980,p8981,p8982,p8983,p8984,p8985,p8986,p8987,p8988,p8989,p8990,p8991,p8992,p8993,p8994,p8995,p8996,p8997,p8998,p8999,p9000,p9001,p9002,p9003,p9004,p9005,p9006,p9007,p9008,p9009,p9010,p9011,p9012,p9013,p9014,p9015,p9016,p9017,p9018,p9019,p9020,p9021,p9022,p9023,p9024,p9025,p9026,p9027,p9028,p9029,p9030,p9031,p9032,p9033,p9034,p9035,p9036,p9037,p9038,p9039,p9040,p9041,p9042,p9043,p9044,p9045,p9046,p9047,p9048,p9049,p9050,p9051,p9052,p9053,p9054,p9055,p9056,p9057,p9058,p9059,p9060,p9061,p9062,p9063,p9064,p9065,p9066,p9067,p9068,p9069,p9070,p9071,p9072,p9073,p9074,p9075,p9076,p9077,p9078,p9079,p9080,p9081,p9082,p9083,p9084,p9085,p9086,p9087,p9088,p9089,p9090,p9091,p9092,p9093,p9094,p9095,p9096,p9097,p9098,p9099,p9100,p9101,p9102,p9103,p9104,p9105,p9106,p9107,p9108,p9109,p9110,p9111,p9112,p9113,p9114,p9115,p9116,p9117,p9118,p9119,p9120,p9121,p9122,p9123,p9124,p9125,p9126,p9127,p9128,p9129,p9130,p9131,p9132,p9133,p9134,p9135,p9136,p9137,p9138,p9139,p9140,p9141,p9142,p9143,p9144,p9145,p9146,p9147,p9148,p9149,p9150,p9151,p9152,p9153,p9154,p9155,p9156,p9157,p9158,p9159,p9160,p9161,p9162,p9163,p9164,p9165,p9166,p9167,p9168,p9169,p9170,p9171,p9172,p9173,p9174,p9175,p9176,p9177,p9178,p9179,p9180,p9181,p9182,p9183,p9184,p9185,p9186,p9187,p9188,p9189,p9190,p9191,p9192,p9193,p9194,p9195,p9196,p9197,p9198,p9199,p9200,p9201,p9202,p9203,p9204,p9205,p9206,p9207,p9208,p9209,p9210,p9211,p9212,p9213,p9214,p9215,p9216,p9217,p9218,p9219,p9220,p9221,p9222,p9223,p9224,p9225,p9226,p9227,p9228,p9229,p9230,p9231,p9232,p9233,p9234,p9235,p9236,p9237,p9238,p9239,p9240,p9241,p9242,p9243,p9244,p9245,p9246,p9247,p9248,p9249,p9250,p9251,p9252,p9253,p9254,p9255,p9256,p9257,p9258,p9259,p9260,p9261,p9262,p9263,p9264,p9265,p9266,p9267,p9268,p9269,p9270,p9271,p9272,p9273,p9274,p9275,p9276,p9277,p9278,p9279,p9280,p9281,p9282,p9283,p9284,p9285,p9286,p9287,p9288,p9289,p9290,p9291,p9292,p9293,p9294,p9295,p9296,p9297,p9298,p9299,p9300,p9301,p9302,p9303,p9304,p9305,p9306,p9307,p9308,p9309,p9310,p9311,p9312,p9313,p9314,p9315,p9316,p9317,p9318,p9319,p9320,p9321,p9322,p9323,p9324,p9325,p9326,p9327,p9328,p9329,p9330,p9331,p9332,p9333,p9334,p9335,p9336,p9337,p9338,p9339,p9340,p9341,p9342,p9343,p9344,p9345,p9346,p9347,p9348,p9349,p9350,p9351,p9352,p9353,p9354,p9355,p9356,p9357,p9358,p9359,p9360,p9361,p9362,p9363,p9364,p9365,p9366,p9367,p9368,p9369,p9370,p9371,p9372,p9373,p9374,p9375,p9376,p9377,p9378,p9379,p9380,p9381,p9382,p9383,p9384,p9385,p9386,p9387,p9388,p9389,p9390,p9391,p9392,p9393,p9394,p9395,p9396,p9397,p9398,p9399,p9400,p9401,p9402,p9403,p9404,p9405,p9406,p9407,p9408,p9409,p9410,p9411,p9412,p9413,p9414,p9415,p9416,p9417,p9418,p9419,p9420,p9421,p9422,p9423,p9424,p9425,p9426,p9427,p9428,p9429,p9430,p9431,p9432,p9433,p9434,p9435,p9436,p9437,p9438,p9439,p9440,p9441,p9442,p9443,p9444,p9445,p9446,p9447,p9448,p9449,p9450,p9451,p9452,p9453,p9454,p9455,p9456,p9457,p9458,p9459,p9460,p9461,p9462,p9463,p9464,p9465,p9466,p9467,p9468,p9469,p9470,p9471,p9472,p9473,p9474,p9475,p9476,p9477,p9478,p9479,p9480,p9481,p9482,p9483,p9484,p9485,p9486,p9487,p9488,p9489,p9490,p9491,p9492,p9493,p9494,p9495,p9496,p9497,p9498,p9499,p9500,p9501,p9502,p9503,p9504,p9505,p9506,p9507,p9508,p9509,p9510,p9511,p9512,p9513,p9514,p9515,p9516,p9517,p9518,p9519,p9520,p9521,p9522,p9523,p9524,p9525,p9526,p9527,p9528,p9529,p9530,p9531,p9532,p9533,p9534,p9535,p9536,p9537,p9538,p9539,p9540,p9541,p9542,p9543,p9544,p9545,p9546,p9547,p9548,p9549,p9550,p9551,p9552,p9553,p9554,p9555,p9556,p9557,p9558,p9559,p9560,p9561,p9562,p9563,p9564,p9565,p9566,p9567,p9568,p9569,p9570,p9571,p9572,p9573,p9574,p9575,p9576,p9577,p9578,p9579,p9580,p9581,p9582,p9583,p9584,p9585,p9586,p9587,p9588,p9589,p9590,p9591,p9592,p9593,p9594,p9595,p9596,p9597,p9598,p9599,p9600,p9601,p9602,p9603,p9604,p9605,p9606,p9607,p9608,p9609,p9610,p9611,p9612,p9613,p9614,p9615,p9616,p9617,p9618,p9619,p9620,p9621,p9622,p9623,p9624,p9625,p9626,p9627,p9628,p9629,p9630,p9631,p9632,p9633,p9634,p9635,p9636,p9637,p9638,p9639,p9640,p9641,p9642,p9643,p9644,p9645,p9646,p9647,p9648,p9649,p9650,p9651,p9652,p9653,p9654,p9655,p9656,p9657,p9658,p9659,p9660,p9661,p9662,p9663,p9664,p9665,p9666,p9667,p9668,p9669,p9670,p9671,p9672,p9673,p9674,p9675,p9676,p9677,p9678,p9679,p9680,p9681,p9682,p9683,p9684,p9685,p9686,p9687,p9688,p9689,p9690,p9691,p9692,p9693,p9694,p9695,p9696,p9697,p9698,p9699,p9700,p9701,p9702,p9703,p9704,p9705;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_0_16,x[0],y[16]);
and and17(ip_0_17,x[0],y[17]);
and and18(ip_0_18,x[0],y[18]);
and and19(ip_0_19,x[0],y[19]);
and and20(ip_0_20,x[0],y[20]);
and and21(ip_0_21,x[0],y[21]);
and and22(ip_0_22,x[0],y[22]);
and and23(ip_0_23,x[0],y[23]);
and and24(ip_0_24,x[0],y[24]);
and and25(ip_0_25,x[0],y[25]);
and and26(ip_0_26,x[0],y[26]);
and and27(ip_0_27,x[0],y[27]);
and and28(ip_0_28,x[0],y[28]);
and and29(ip_0_29,x[0],y[29]);
and and30(ip_0_30,x[0],y[30]);
and and31(ip_0_31,x[0],y[31]);
and and32(ip_0_32,x[0],y[32]);
and and33(ip_0_33,x[0],y[33]);
and and34(ip_0_34,x[0],y[34]);
and and35(ip_0_35,x[0],y[35]);
and and36(ip_0_36,x[0],y[36]);
and and37(ip_0_37,x[0],y[37]);
and and38(ip_0_38,x[0],y[38]);
and and39(ip_0_39,x[0],y[39]);
and and40(ip_0_40,x[0],y[40]);
and and41(ip_0_41,x[0],y[41]);
and and42(ip_0_42,x[0],y[42]);
and and43(ip_0_43,x[0],y[43]);
and and44(ip_0_44,x[0],y[44]);
and and45(ip_0_45,x[0],y[45]);
and and46(ip_0_46,x[0],y[46]);
and and47(ip_0_47,x[0],y[47]);
and and48(ip_0_48,x[0],y[48]);
and and49(ip_0_49,x[0],y[49]);
and and50(ip_0_50,x[0],y[50]);
and and51(ip_0_51,x[0],y[51]);
and and52(ip_0_52,x[0],y[52]);
and and53(ip_0_53,x[0],y[53]);
and and54(ip_0_54,x[0],y[54]);
and and55(ip_0_55,x[0],y[55]);
and and56(ip_0_56,x[0],y[56]);
and and57(ip_0_57,x[0],y[57]);
and and58(ip_0_58,x[0],y[58]);
and and59(ip_0_59,x[0],y[59]);
and and60(ip_0_60,x[0],y[60]);
and and61(ip_0_61,x[0],y[61]);
and and62(ip_0_62,x[0],y[62]);
and and63(ip_0_63,x[0],y[63]);
and and64(ip_1_0,x[1],y[0]);
and and65(ip_1_1,x[1],y[1]);
and and66(ip_1_2,x[1],y[2]);
and and67(ip_1_3,x[1],y[3]);
and and68(ip_1_4,x[1],y[4]);
and and69(ip_1_5,x[1],y[5]);
and and70(ip_1_6,x[1],y[6]);
and and71(ip_1_7,x[1],y[7]);
and and72(ip_1_8,x[1],y[8]);
and and73(ip_1_9,x[1],y[9]);
and and74(ip_1_10,x[1],y[10]);
and and75(ip_1_11,x[1],y[11]);
and and76(ip_1_12,x[1],y[12]);
and and77(ip_1_13,x[1],y[13]);
and and78(ip_1_14,x[1],y[14]);
and and79(ip_1_15,x[1],y[15]);
and and80(ip_1_16,x[1],y[16]);
and and81(ip_1_17,x[1],y[17]);
and and82(ip_1_18,x[1],y[18]);
and and83(ip_1_19,x[1],y[19]);
and and84(ip_1_20,x[1],y[20]);
and and85(ip_1_21,x[1],y[21]);
and and86(ip_1_22,x[1],y[22]);
and and87(ip_1_23,x[1],y[23]);
and and88(ip_1_24,x[1],y[24]);
and and89(ip_1_25,x[1],y[25]);
and and90(ip_1_26,x[1],y[26]);
and and91(ip_1_27,x[1],y[27]);
and and92(ip_1_28,x[1],y[28]);
and and93(ip_1_29,x[1],y[29]);
and and94(ip_1_30,x[1],y[30]);
and and95(ip_1_31,x[1],y[31]);
and and96(ip_1_32,x[1],y[32]);
and and97(ip_1_33,x[1],y[33]);
and and98(ip_1_34,x[1],y[34]);
and and99(ip_1_35,x[1],y[35]);
and and100(ip_1_36,x[1],y[36]);
and and101(ip_1_37,x[1],y[37]);
and and102(ip_1_38,x[1],y[38]);
and and103(ip_1_39,x[1],y[39]);
and and104(ip_1_40,x[1],y[40]);
and and105(ip_1_41,x[1],y[41]);
and and106(ip_1_42,x[1],y[42]);
and and107(ip_1_43,x[1],y[43]);
and and108(ip_1_44,x[1],y[44]);
and and109(ip_1_45,x[1],y[45]);
and and110(ip_1_46,x[1],y[46]);
and and111(ip_1_47,x[1],y[47]);
and and112(ip_1_48,x[1],y[48]);
and and113(ip_1_49,x[1],y[49]);
and and114(ip_1_50,x[1],y[50]);
and and115(ip_1_51,x[1],y[51]);
and and116(ip_1_52,x[1],y[52]);
and and117(ip_1_53,x[1],y[53]);
and and118(ip_1_54,x[1],y[54]);
and and119(ip_1_55,x[1],y[55]);
and and120(ip_1_56,x[1],y[56]);
and and121(ip_1_57,x[1],y[57]);
and and122(ip_1_58,x[1],y[58]);
and and123(ip_1_59,x[1],y[59]);
and and124(ip_1_60,x[1],y[60]);
and and125(ip_1_61,x[1],y[61]);
and and126(ip_1_62,x[1],y[62]);
and and127(ip_1_63,x[1],y[63]);
and and128(ip_2_0,x[2],y[0]);
and and129(ip_2_1,x[2],y[1]);
and and130(ip_2_2,x[2],y[2]);
and and131(ip_2_3,x[2],y[3]);
and and132(ip_2_4,x[2],y[4]);
and and133(ip_2_5,x[2],y[5]);
and and134(ip_2_6,x[2],y[6]);
and and135(ip_2_7,x[2],y[7]);
and and136(ip_2_8,x[2],y[8]);
and and137(ip_2_9,x[2],y[9]);
and and138(ip_2_10,x[2],y[10]);
and and139(ip_2_11,x[2],y[11]);
and and140(ip_2_12,x[2],y[12]);
and and141(ip_2_13,x[2],y[13]);
and and142(ip_2_14,x[2],y[14]);
and and143(ip_2_15,x[2],y[15]);
and and144(ip_2_16,x[2],y[16]);
and and145(ip_2_17,x[2],y[17]);
and and146(ip_2_18,x[2],y[18]);
and and147(ip_2_19,x[2],y[19]);
and and148(ip_2_20,x[2],y[20]);
and and149(ip_2_21,x[2],y[21]);
and and150(ip_2_22,x[2],y[22]);
and and151(ip_2_23,x[2],y[23]);
and and152(ip_2_24,x[2],y[24]);
and and153(ip_2_25,x[2],y[25]);
and and154(ip_2_26,x[2],y[26]);
and and155(ip_2_27,x[2],y[27]);
and and156(ip_2_28,x[2],y[28]);
and and157(ip_2_29,x[2],y[29]);
and and158(ip_2_30,x[2],y[30]);
and and159(ip_2_31,x[2],y[31]);
and and160(ip_2_32,x[2],y[32]);
and and161(ip_2_33,x[2],y[33]);
and and162(ip_2_34,x[2],y[34]);
and and163(ip_2_35,x[2],y[35]);
and and164(ip_2_36,x[2],y[36]);
and and165(ip_2_37,x[2],y[37]);
and and166(ip_2_38,x[2],y[38]);
and and167(ip_2_39,x[2],y[39]);
and and168(ip_2_40,x[2],y[40]);
and and169(ip_2_41,x[2],y[41]);
and and170(ip_2_42,x[2],y[42]);
and and171(ip_2_43,x[2],y[43]);
and and172(ip_2_44,x[2],y[44]);
and and173(ip_2_45,x[2],y[45]);
and and174(ip_2_46,x[2],y[46]);
and and175(ip_2_47,x[2],y[47]);
and and176(ip_2_48,x[2],y[48]);
and and177(ip_2_49,x[2],y[49]);
and and178(ip_2_50,x[2],y[50]);
and and179(ip_2_51,x[2],y[51]);
and and180(ip_2_52,x[2],y[52]);
and and181(ip_2_53,x[2],y[53]);
and and182(ip_2_54,x[2],y[54]);
and and183(ip_2_55,x[2],y[55]);
and and184(ip_2_56,x[2],y[56]);
and and185(ip_2_57,x[2],y[57]);
and and186(ip_2_58,x[2],y[58]);
and and187(ip_2_59,x[2],y[59]);
and and188(ip_2_60,x[2],y[60]);
and and189(ip_2_61,x[2],y[61]);
and and190(ip_2_62,x[2],y[62]);
and and191(ip_2_63,x[2],y[63]);
and and192(ip_3_0,x[3],y[0]);
and and193(ip_3_1,x[3],y[1]);
and and194(ip_3_2,x[3],y[2]);
and and195(ip_3_3,x[3],y[3]);
and and196(ip_3_4,x[3],y[4]);
and and197(ip_3_5,x[3],y[5]);
and and198(ip_3_6,x[3],y[6]);
and and199(ip_3_7,x[3],y[7]);
and and200(ip_3_8,x[3],y[8]);
and and201(ip_3_9,x[3],y[9]);
and and202(ip_3_10,x[3],y[10]);
and and203(ip_3_11,x[3],y[11]);
and and204(ip_3_12,x[3],y[12]);
and and205(ip_3_13,x[3],y[13]);
and and206(ip_3_14,x[3],y[14]);
and and207(ip_3_15,x[3],y[15]);
and and208(ip_3_16,x[3],y[16]);
and and209(ip_3_17,x[3],y[17]);
and and210(ip_3_18,x[3],y[18]);
and and211(ip_3_19,x[3],y[19]);
and and212(ip_3_20,x[3],y[20]);
and and213(ip_3_21,x[3],y[21]);
and and214(ip_3_22,x[3],y[22]);
and and215(ip_3_23,x[3],y[23]);
and and216(ip_3_24,x[3],y[24]);
and and217(ip_3_25,x[3],y[25]);
and and218(ip_3_26,x[3],y[26]);
and and219(ip_3_27,x[3],y[27]);
and and220(ip_3_28,x[3],y[28]);
and and221(ip_3_29,x[3],y[29]);
and and222(ip_3_30,x[3],y[30]);
and and223(ip_3_31,x[3],y[31]);
and and224(ip_3_32,x[3],y[32]);
and and225(ip_3_33,x[3],y[33]);
and and226(ip_3_34,x[3],y[34]);
and and227(ip_3_35,x[3],y[35]);
and and228(ip_3_36,x[3],y[36]);
and and229(ip_3_37,x[3],y[37]);
and and230(ip_3_38,x[3],y[38]);
and and231(ip_3_39,x[3],y[39]);
and and232(ip_3_40,x[3],y[40]);
and and233(ip_3_41,x[3],y[41]);
and and234(ip_3_42,x[3],y[42]);
and and235(ip_3_43,x[3],y[43]);
and and236(ip_3_44,x[3],y[44]);
and and237(ip_3_45,x[3],y[45]);
and and238(ip_3_46,x[3],y[46]);
and and239(ip_3_47,x[3],y[47]);
and and240(ip_3_48,x[3],y[48]);
and and241(ip_3_49,x[3],y[49]);
and and242(ip_3_50,x[3],y[50]);
and and243(ip_3_51,x[3],y[51]);
and and244(ip_3_52,x[3],y[52]);
and and245(ip_3_53,x[3],y[53]);
and and246(ip_3_54,x[3],y[54]);
and and247(ip_3_55,x[3],y[55]);
and and248(ip_3_56,x[3],y[56]);
and and249(ip_3_57,x[3],y[57]);
and and250(ip_3_58,x[3],y[58]);
and and251(ip_3_59,x[3],y[59]);
and and252(ip_3_60,x[3],y[60]);
and and253(ip_3_61,x[3],y[61]);
and and254(ip_3_62,x[3],y[62]);
and and255(ip_3_63,x[3],y[63]);
and and256(ip_4_0,x[4],y[0]);
and and257(ip_4_1,x[4],y[1]);
and and258(ip_4_2,x[4],y[2]);
and and259(ip_4_3,x[4],y[3]);
and and260(ip_4_4,x[4],y[4]);
and and261(ip_4_5,x[4],y[5]);
and and262(ip_4_6,x[4],y[6]);
and and263(ip_4_7,x[4],y[7]);
and and264(ip_4_8,x[4],y[8]);
and and265(ip_4_9,x[4],y[9]);
and and266(ip_4_10,x[4],y[10]);
and and267(ip_4_11,x[4],y[11]);
and and268(ip_4_12,x[4],y[12]);
and and269(ip_4_13,x[4],y[13]);
and and270(ip_4_14,x[4],y[14]);
and and271(ip_4_15,x[4],y[15]);
and and272(ip_4_16,x[4],y[16]);
and and273(ip_4_17,x[4],y[17]);
and and274(ip_4_18,x[4],y[18]);
and and275(ip_4_19,x[4],y[19]);
and and276(ip_4_20,x[4],y[20]);
and and277(ip_4_21,x[4],y[21]);
and and278(ip_4_22,x[4],y[22]);
and and279(ip_4_23,x[4],y[23]);
and and280(ip_4_24,x[4],y[24]);
and and281(ip_4_25,x[4],y[25]);
and and282(ip_4_26,x[4],y[26]);
and and283(ip_4_27,x[4],y[27]);
and and284(ip_4_28,x[4],y[28]);
and and285(ip_4_29,x[4],y[29]);
and and286(ip_4_30,x[4],y[30]);
and and287(ip_4_31,x[4],y[31]);
and and288(ip_4_32,x[4],y[32]);
and and289(ip_4_33,x[4],y[33]);
and and290(ip_4_34,x[4],y[34]);
and and291(ip_4_35,x[4],y[35]);
and and292(ip_4_36,x[4],y[36]);
and and293(ip_4_37,x[4],y[37]);
and and294(ip_4_38,x[4],y[38]);
and and295(ip_4_39,x[4],y[39]);
and and296(ip_4_40,x[4],y[40]);
and and297(ip_4_41,x[4],y[41]);
and and298(ip_4_42,x[4],y[42]);
and and299(ip_4_43,x[4],y[43]);
and and300(ip_4_44,x[4],y[44]);
and and301(ip_4_45,x[4],y[45]);
and and302(ip_4_46,x[4],y[46]);
and and303(ip_4_47,x[4],y[47]);
and and304(ip_4_48,x[4],y[48]);
and and305(ip_4_49,x[4],y[49]);
and and306(ip_4_50,x[4],y[50]);
and and307(ip_4_51,x[4],y[51]);
and and308(ip_4_52,x[4],y[52]);
and and309(ip_4_53,x[4],y[53]);
and and310(ip_4_54,x[4],y[54]);
and and311(ip_4_55,x[4],y[55]);
and and312(ip_4_56,x[4],y[56]);
and and313(ip_4_57,x[4],y[57]);
and and314(ip_4_58,x[4],y[58]);
and and315(ip_4_59,x[4],y[59]);
and and316(ip_4_60,x[4],y[60]);
and and317(ip_4_61,x[4],y[61]);
and and318(ip_4_62,x[4],y[62]);
and and319(ip_4_63,x[4],y[63]);
and and320(ip_5_0,x[5],y[0]);
and and321(ip_5_1,x[5],y[1]);
and and322(ip_5_2,x[5],y[2]);
and and323(ip_5_3,x[5],y[3]);
and and324(ip_5_4,x[5],y[4]);
and and325(ip_5_5,x[5],y[5]);
and and326(ip_5_6,x[5],y[6]);
and and327(ip_5_7,x[5],y[7]);
and and328(ip_5_8,x[5],y[8]);
and and329(ip_5_9,x[5],y[9]);
and and330(ip_5_10,x[5],y[10]);
and and331(ip_5_11,x[5],y[11]);
and and332(ip_5_12,x[5],y[12]);
and and333(ip_5_13,x[5],y[13]);
and and334(ip_5_14,x[5],y[14]);
and and335(ip_5_15,x[5],y[15]);
and and336(ip_5_16,x[5],y[16]);
and and337(ip_5_17,x[5],y[17]);
and and338(ip_5_18,x[5],y[18]);
and and339(ip_5_19,x[5],y[19]);
and and340(ip_5_20,x[5],y[20]);
and and341(ip_5_21,x[5],y[21]);
and and342(ip_5_22,x[5],y[22]);
and and343(ip_5_23,x[5],y[23]);
and and344(ip_5_24,x[5],y[24]);
and and345(ip_5_25,x[5],y[25]);
and and346(ip_5_26,x[5],y[26]);
and and347(ip_5_27,x[5],y[27]);
and and348(ip_5_28,x[5],y[28]);
and and349(ip_5_29,x[5],y[29]);
and and350(ip_5_30,x[5],y[30]);
and and351(ip_5_31,x[5],y[31]);
and and352(ip_5_32,x[5],y[32]);
and and353(ip_5_33,x[5],y[33]);
and and354(ip_5_34,x[5],y[34]);
and and355(ip_5_35,x[5],y[35]);
and and356(ip_5_36,x[5],y[36]);
and and357(ip_5_37,x[5],y[37]);
and and358(ip_5_38,x[5],y[38]);
and and359(ip_5_39,x[5],y[39]);
and and360(ip_5_40,x[5],y[40]);
and and361(ip_5_41,x[5],y[41]);
and and362(ip_5_42,x[5],y[42]);
and and363(ip_5_43,x[5],y[43]);
and and364(ip_5_44,x[5],y[44]);
and and365(ip_5_45,x[5],y[45]);
and and366(ip_5_46,x[5],y[46]);
and and367(ip_5_47,x[5],y[47]);
and and368(ip_5_48,x[5],y[48]);
and and369(ip_5_49,x[5],y[49]);
and and370(ip_5_50,x[5],y[50]);
and and371(ip_5_51,x[5],y[51]);
and and372(ip_5_52,x[5],y[52]);
and and373(ip_5_53,x[5],y[53]);
and and374(ip_5_54,x[5],y[54]);
and and375(ip_5_55,x[5],y[55]);
and and376(ip_5_56,x[5],y[56]);
and and377(ip_5_57,x[5],y[57]);
and and378(ip_5_58,x[5],y[58]);
and and379(ip_5_59,x[5],y[59]);
and and380(ip_5_60,x[5],y[60]);
and and381(ip_5_61,x[5],y[61]);
and and382(ip_5_62,x[5],y[62]);
and and383(ip_5_63,x[5],y[63]);
and and384(ip_6_0,x[6],y[0]);
and and385(ip_6_1,x[6],y[1]);
and and386(ip_6_2,x[6],y[2]);
and and387(ip_6_3,x[6],y[3]);
and and388(ip_6_4,x[6],y[4]);
and and389(ip_6_5,x[6],y[5]);
and and390(ip_6_6,x[6],y[6]);
and and391(ip_6_7,x[6],y[7]);
and and392(ip_6_8,x[6],y[8]);
and and393(ip_6_9,x[6],y[9]);
and and394(ip_6_10,x[6],y[10]);
and and395(ip_6_11,x[6],y[11]);
and and396(ip_6_12,x[6],y[12]);
and and397(ip_6_13,x[6],y[13]);
and and398(ip_6_14,x[6],y[14]);
and and399(ip_6_15,x[6],y[15]);
and and400(ip_6_16,x[6],y[16]);
and and401(ip_6_17,x[6],y[17]);
and and402(ip_6_18,x[6],y[18]);
and and403(ip_6_19,x[6],y[19]);
and and404(ip_6_20,x[6],y[20]);
and and405(ip_6_21,x[6],y[21]);
and and406(ip_6_22,x[6],y[22]);
and and407(ip_6_23,x[6],y[23]);
and and408(ip_6_24,x[6],y[24]);
and and409(ip_6_25,x[6],y[25]);
and and410(ip_6_26,x[6],y[26]);
and and411(ip_6_27,x[6],y[27]);
and and412(ip_6_28,x[6],y[28]);
and and413(ip_6_29,x[6],y[29]);
and and414(ip_6_30,x[6],y[30]);
and and415(ip_6_31,x[6],y[31]);
and and416(ip_6_32,x[6],y[32]);
and and417(ip_6_33,x[6],y[33]);
and and418(ip_6_34,x[6],y[34]);
and and419(ip_6_35,x[6],y[35]);
and and420(ip_6_36,x[6],y[36]);
and and421(ip_6_37,x[6],y[37]);
and and422(ip_6_38,x[6],y[38]);
and and423(ip_6_39,x[6],y[39]);
and and424(ip_6_40,x[6],y[40]);
and and425(ip_6_41,x[6],y[41]);
and and426(ip_6_42,x[6],y[42]);
and and427(ip_6_43,x[6],y[43]);
and and428(ip_6_44,x[6],y[44]);
and and429(ip_6_45,x[6],y[45]);
and and430(ip_6_46,x[6],y[46]);
and and431(ip_6_47,x[6],y[47]);
and and432(ip_6_48,x[6],y[48]);
and and433(ip_6_49,x[6],y[49]);
and and434(ip_6_50,x[6],y[50]);
and and435(ip_6_51,x[6],y[51]);
and and436(ip_6_52,x[6],y[52]);
and and437(ip_6_53,x[6],y[53]);
and and438(ip_6_54,x[6],y[54]);
and and439(ip_6_55,x[6],y[55]);
and and440(ip_6_56,x[6],y[56]);
and and441(ip_6_57,x[6],y[57]);
and and442(ip_6_58,x[6],y[58]);
and and443(ip_6_59,x[6],y[59]);
and and444(ip_6_60,x[6],y[60]);
and and445(ip_6_61,x[6],y[61]);
and and446(ip_6_62,x[6],y[62]);
and and447(ip_6_63,x[6],y[63]);
and and448(ip_7_0,x[7],y[0]);
and and449(ip_7_1,x[7],y[1]);
and and450(ip_7_2,x[7],y[2]);
and and451(ip_7_3,x[7],y[3]);
and and452(ip_7_4,x[7],y[4]);
and and453(ip_7_5,x[7],y[5]);
and and454(ip_7_6,x[7],y[6]);
and and455(ip_7_7,x[7],y[7]);
and and456(ip_7_8,x[7],y[8]);
and and457(ip_7_9,x[7],y[9]);
and and458(ip_7_10,x[7],y[10]);
and and459(ip_7_11,x[7],y[11]);
and and460(ip_7_12,x[7],y[12]);
and and461(ip_7_13,x[7],y[13]);
and and462(ip_7_14,x[7],y[14]);
and and463(ip_7_15,x[7],y[15]);
and and464(ip_7_16,x[7],y[16]);
and and465(ip_7_17,x[7],y[17]);
and and466(ip_7_18,x[7],y[18]);
and and467(ip_7_19,x[7],y[19]);
and and468(ip_7_20,x[7],y[20]);
and and469(ip_7_21,x[7],y[21]);
and and470(ip_7_22,x[7],y[22]);
and and471(ip_7_23,x[7],y[23]);
and and472(ip_7_24,x[7],y[24]);
and and473(ip_7_25,x[7],y[25]);
and and474(ip_7_26,x[7],y[26]);
and and475(ip_7_27,x[7],y[27]);
and and476(ip_7_28,x[7],y[28]);
and and477(ip_7_29,x[7],y[29]);
and and478(ip_7_30,x[7],y[30]);
and and479(ip_7_31,x[7],y[31]);
and and480(ip_7_32,x[7],y[32]);
and and481(ip_7_33,x[7],y[33]);
and and482(ip_7_34,x[7],y[34]);
and and483(ip_7_35,x[7],y[35]);
and and484(ip_7_36,x[7],y[36]);
and and485(ip_7_37,x[7],y[37]);
and and486(ip_7_38,x[7],y[38]);
and and487(ip_7_39,x[7],y[39]);
and and488(ip_7_40,x[7],y[40]);
and and489(ip_7_41,x[7],y[41]);
and and490(ip_7_42,x[7],y[42]);
and and491(ip_7_43,x[7],y[43]);
and and492(ip_7_44,x[7],y[44]);
and and493(ip_7_45,x[7],y[45]);
and and494(ip_7_46,x[7],y[46]);
and and495(ip_7_47,x[7],y[47]);
and and496(ip_7_48,x[7],y[48]);
and and497(ip_7_49,x[7],y[49]);
and and498(ip_7_50,x[7],y[50]);
and and499(ip_7_51,x[7],y[51]);
and and500(ip_7_52,x[7],y[52]);
and and501(ip_7_53,x[7],y[53]);
and and502(ip_7_54,x[7],y[54]);
and and503(ip_7_55,x[7],y[55]);
and and504(ip_7_56,x[7],y[56]);
and and505(ip_7_57,x[7],y[57]);
and and506(ip_7_58,x[7],y[58]);
and and507(ip_7_59,x[7],y[59]);
and and508(ip_7_60,x[7],y[60]);
and and509(ip_7_61,x[7],y[61]);
and and510(ip_7_62,x[7],y[62]);
and and511(ip_7_63,x[7],y[63]);
and and512(ip_8_0,x[8],y[0]);
and and513(ip_8_1,x[8],y[1]);
and and514(ip_8_2,x[8],y[2]);
and and515(ip_8_3,x[8],y[3]);
and and516(ip_8_4,x[8],y[4]);
and and517(ip_8_5,x[8],y[5]);
and and518(ip_8_6,x[8],y[6]);
and and519(ip_8_7,x[8],y[7]);
and and520(ip_8_8,x[8],y[8]);
and and521(ip_8_9,x[8],y[9]);
and and522(ip_8_10,x[8],y[10]);
and and523(ip_8_11,x[8],y[11]);
and and524(ip_8_12,x[8],y[12]);
and and525(ip_8_13,x[8],y[13]);
and and526(ip_8_14,x[8],y[14]);
and and527(ip_8_15,x[8],y[15]);
and and528(ip_8_16,x[8],y[16]);
and and529(ip_8_17,x[8],y[17]);
and and530(ip_8_18,x[8],y[18]);
and and531(ip_8_19,x[8],y[19]);
and and532(ip_8_20,x[8],y[20]);
and and533(ip_8_21,x[8],y[21]);
and and534(ip_8_22,x[8],y[22]);
and and535(ip_8_23,x[8],y[23]);
and and536(ip_8_24,x[8],y[24]);
and and537(ip_8_25,x[8],y[25]);
and and538(ip_8_26,x[8],y[26]);
and and539(ip_8_27,x[8],y[27]);
and and540(ip_8_28,x[8],y[28]);
and and541(ip_8_29,x[8],y[29]);
and and542(ip_8_30,x[8],y[30]);
and and543(ip_8_31,x[8],y[31]);
and and544(ip_8_32,x[8],y[32]);
and and545(ip_8_33,x[8],y[33]);
and and546(ip_8_34,x[8],y[34]);
and and547(ip_8_35,x[8],y[35]);
and and548(ip_8_36,x[8],y[36]);
and and549(ip_8_37,x[8],y[37]);
and and550(ip_8_38,x[8],y[38]);
and and551(ip_8_39,x[8],y[39]);
and and552(ip_8_40,x[8],y[40]);
and and553(ip_8_41,x[8],y[41]);
and and554(ip_8_42,x[8],y[42]);
and and555(ip_8_43,x[8],y[43]);
and and556(ip_8_44,x[8],y[44]);
and and557(ip_8_45,x[8],y[45]);
and and558(ip_8_46,x[8],y[46]);
and and559(ip_8_47,x[8],y[47]);
and and560(ip_8_48,x[8],y[48]);
and and561(ip_8_49,x[8],y[49]);
and and562(ip_8_50,x[8],y[50]);
and and563(ip_8_51,x[8],y[51]);
and and564(ip_8_52,x[8],y[52]);
and and565(ip_8_53,x[8],y[53]);
and and566(ip_8_54,x[8],y[54]);
and and567(ip_8_55,x[8],y[55]);
and and568(ip_8_56,x[8],y[56]);
and and569(ip_8_57,x[8],y[57]);
and and570(ip_8_58,x[8],y[58]);
and and571(ip_8_59,x[8],y[59]);
and and572(ip_8_60,x[8],y[60]);
and and573(ip_8_61,x[8],y[61]);
and and574(ip_8_62,x[8],y[62]);
and and575(ip_8_63,x[8],y[63]);
and and576(ip_9_0,x[9],y[0]);
and and577(ip_9_1,x[9],y[1]);
and and578(ip_9_2,x[9],y[2]);
and and579(ip_9_3,x[9],y[3]);
and and580(ip_9_4,x[9],y[4]);
and and581(ip_9_5,x[9],y[5]);
and and582(ip_9_6,x[9],y[6]);
and and583(ip_9_7,x[9],y[7]);
and and584(ip_9_8,x[9],y[8]);
and and585(ip_9_9,x[9],y[9]);
and and586(ip_9_10,x[9],y[10]);
and and587(ip_9_11,x[9],y[11]);
and and588(ip_9_12,x[9],y[12]);
and and589(ip_9_13,x[9],y[13]);
and and590(ip_9_14,x[9],y[14]);
and and591(ip_9_15,x[9],y[15]);
and and592(ip_9_16,x[9],y[16]);
and and593(ip_9_17,x[9],y[17]);
and and594(ip_9_18,x[9],y[18]);
and and595(ip_9_19,x[9],y[19]);
and and596(ip_9_20,x[9],y[20]);
and and597(ip_9_21,x[9],y[21]);
and and598(ip_9_22,x[9],y[22]);
and and599(ip_9_23,x[9],y[23]);
and and600(ip_9_24,x[9],y[24]);
and and601(ip_9_25,x[9],y[25]);
and and602(ip_9_26,x[9],y[26]);
and and603(ip_9_27,x[9],y[27]);
and and604(ip_9_28,x[9],y[28]);
and and605(ip_9_29,x[9],y[29]);
and and606(ip_9_30,x[9],y[30]);
and and607(ip_9_31,x[9],y[31]);
and and608(ip_9_32,x[9],y[32]);
and and609(ip_9_33,x[9],y[33]);
and and610(ip_9_34,x[9],y[34]);
and and611(ip_9_35,x[9],y[35]);
and and612(ip_9_36,x[9],y[36]);
and and613(ip_9_37,x[9],y[37]);
and and614(ip_9_38,x[9],y[38]);
and and615(ip_9_39,x[9],y[39]);
and and616(ip_9_40,x[9],y[40]);
and and617(ip_9_41,x[9],y[41]);
and and618(ip_9_42,x[9],y[42]);
and and619(ip_9_43,x[9],y[43]);
and and620(ip_9_44,x[9],y[44]);
and and621(ip_9_45,x[9],y[45]);
and and622(ip_9_46,x[9],y[46]);
and and623(ip_9_47,x[9],y[47]);
and and624(ip_9_48,x[9],y[48]);
and and625(ip_9_49,x[9],y[49]);
and and626(ip_9_50,x[9],y[50]);
and and627(ip_9_51,x[9],y[51]);
and and628(ip_9_52,x[9],y[52]);
and and629(ip_9_53,x[9],y[53]);
and and630(ip_9_54,x[9],y[54]);
and and631(ip_9_55,x[9],y[55]);
and and632(ip_9_56,x[9],y[56]);
and and633(ip_9_57,x[9],y[57]);
and and634(ip_9_58,x[9],y[58]);
and and635(ip_9_59,x[9],y[59]);
and and636(ip_9_60,x[9],y[60]);
and and637(ip_9_61,x[9],y[61]);
and and638(ip_9_62,x[9],y[62]);
and and639(ip_9_63,x[9],y[63]);
and and640(ip_10_0,x[10],y[0]);
and and641(ip_10_1,x[10],y[1]);
and and642(ip_10_2,x[10],y[2]);
and and643(ip_10_3,x[10],y[3]);
and and644(ip_10_4,x[10],y[4]);
and and645(ip_10_5,x[10],y[5]);
and and646(ip_10_6,x[10],y[6]);
and and647(ip_10_7,x[10],y[7]);
and and648(ip_10_8,x[10],y[8]);
and and649(ip_10_9,x[10],y[9]);
and and650(ip_10_10,x[10],y[10]);
and and651(ip_10_11,x[10],y[11]);
and and652(ip_10_12,x[10],y[12]);
and and653(ip_10_13,x[10],y[13]);
and and654(ip_10_14,x[10],y[14]);
and and655(ip_10_15,x[10],y[15]);
and and656(ip_10_16,x[10],y[16]);
and and657(ip_10_17,x[10],y[17]);
and and658(ip_10_18,x[10],y[18]);
and and659(ip_10_19,x[10],y[19]);
and and660(ip_10_20,x[10],y[20]);
and and661(ip_10_21,x[10],y[21]);
and and662(ip_10_22,x[10],y[22]);
and and663(ip_10_23,x[10],y[23]);
and and664(ip_10_24,x[10],y[24]);
and and665(ip_10_25,x[10],y[25]);
and and666(ip_10_26,x[10],y[26]);
and and667(ip_10_27,x[10],y[27]);
and and668(ip_10_28,x[10],y[28]);
and and669(ip_10_29,x[10],y[29]);
and and670(ip_10_30,x[10],y[30]);
and and671(ip_10_31,x[10],y[31]);
and and672(ip_10_32,x[10],y[32]);
and and673(ip_10_33,x[10],y[33]);
and and674(ip_10_34,x[10],y[34]);
and and675(ip_10_35,x[10],y[35]);
and and676(ip_10_36,x[10],y[36]);
and and677(ip_10_37,x[10],y[37]);
and and678(ip_10_38,x[10],y[38]);
and and679(ip_10_39,x[10],y[39]);
and and680(ip_10_40,x[10],y[40]);
and and681(ip_10_41,x[10],y[41]);
and and682(ip_10_42,x[10],y[42]);
and and683(ip_10_43,x[10],y[43]);
and and684(ip_10_44,x[10],y[44]);
and and685(ip_10_45,x[10],y[45]);
and and686(ip_10_46,x[10],y[46]);
and and687(ip_10_47,x[10],y[47]);
and and688(ip_10_48,x[10],y[48]);
and and689(ip_10_49,x[10],y[49]);
and and690(ip_10_50,x[10],y[50]);
and and691(ip_10_51,x[10],y[51]);
and and692(ip_10_52,x[10],y[52]);
and and693(ip_10_53,x[10],y[53]);
and and694(ip_10_54,x[10],y[54]);
and and695(ip_10_55,x[10],y[55]);
and and696(ip_10_56,x[10],y[56]);
and and697(ip_10_57,x[10],y[57]);
and and698(ip_10_58,x[10],y[58]);
and and699(ip_10_59,x[10],y[59]);
and and700(ip_10_60,x[10],y[60]);
and and701(ip_10_61,x[10],y[61]);
and and702(ip_10_62,x[10],y[62]);
and and703(ip_10_63,x[10],y[63]);
and and704(ip_11_0,x[11],y[0]);
and and705(ip_11_1,x[11],y[1]);
and and706(ip_11_2,x[11],y[2]);
and and707(ip_11_3,x[11],y[3]);
and and708(ip_11_4,x[11],y[4]);
and and709(ip_11_5,x[11],y[5]);
and and710(ip_11_6,x[11],y[6]);
and and711(ip_11_7,x[11],y[7]);
and and712(ip_11_8,x[11],y[8]);
and and713(ip_11_9,x[11],y[9]);
and and714(ip_11_10,x[11],y[10]);
and and715(ip_11_11,x[11],y[11]);
and and716(ip_11_12,x[11],y[12]);
and and717(ip_11_13,x[11],y[13]);
and and718(ip_11_14,x[11],y[14]);
and and719(ip_11_15,x[11],y[15]);
and and720(ip_11_16,x[11],y[16]);
and and721(ip_11_17,x[11],y[17]);
and and722(ip_11_18,x[11],y[18]);
and and723(ip_11_19,x[11],y[19]);
and and724(ip_11_20,x[11],y[20]);
and and725(ip_11_21,x[11],y[21]);
and and726(ip_11_22,x[11],y[22]);
and and727(ip_11_23,x[11],y[23]);
and and728(ip_11_24,x[11],y[24]);
and and729(ip_11_25,x[11],y[25]);
and and730(ip_11_26,x[11],y[26]);
and and731(ip_11_27,x[11],y[27]);
and and732(ip_11_28,x[11],y[28]);
and and733(ip_11_29,x[11],y[29]);
and and734(ip_11_30,x[11],y[30]);
and and735(ip_11_31,x[11],y[31]);
and and736(ip_11_32,x[11],y[32]);
and and737(ip_11_33,x[11],y[33]);
and and738(ip_11_34,x[11],y[34]);
and and739(ip_11_35,x[11],y[35]);
and and740(ip_11_36,x[11],y[36]);
and and741(ip_11_37,x[11],y[37]);
and and742(ip_11_38,x[11],y[38]);
and and743(ip_11_39,x[11],y[39]);
and and744(ip_11_40,x[11],y[40]);
and and745(ip_11_41,x[11],y[41]);
and and746(ip_11_42,x[11],y[42]);
and and747(ip_11_43,x[11],y[43]);
and and748(ip_11_44,x[11],y[44]);
and and749(ip_11_45,x[11],y[45]);
and and750(ip_11_46,x[11],y[46]);
and and751(ip_11_47,x[11],y[47]);
and and752(ip_11_48,x[11],y[48]);
and and753(ip_11_49,x[11],y[49]);
and and754(ip_11_50,x[11],y[50]);
and and755(ip_11_51,x[11],y[51]);
and and756(ip_11_52,x[11],y[52]);
and and757(ip_11_53,x[11],y[53]);
and and758(ip_11_54,x[11],y[54]);
and and759(ip_11_55,x[11],y[55]);
and and760(ip_11_56,x[11],y[56]);
and and761(ip_11_57,x[11],y[57]);
and and762(ip_11_58,x[11],y[58]);
and and763(ip_11_59,x[11],y[59]);
and and764(ip_11_60,x[11],y[60]);
and and765(ip_11_61,x[11],y[61]);
and and766(ip_11_62,x[11],y[62]);
and and767(ip_11_63,x[11],y[63]);
and and768(ip_12_0,x[12],y[0]);
and and769(ip_12_1,x[12],y[1]);
and and770(ip_12_2,x[12],y[2]);
and and771(ip_12_3,x[12],y[3]);
and and772(ip_12_4,x[12],y[4]);
and and773(ip_12_5,x[12],y[5]);
and and774(ip_12_6,x[12],y[6]);
and and775(ip_12_7,x[12],y[7]);
and and776(ip_12_8,x[12],y[8]);
and and777(ip_12_9,x[12],y[9]);
and and778(ip_12_10,x[12],y[10]);
and and779(ip_12_11,x[12],y[11]);
and and780(ip_12_12,x[12],y[12]);
and and781(ip_12_13,x[12],y[13]);
and and782(ip_12_14,x[12],y[14]);
and and783(ip_12_15,x[12],y[15]);
and and784(ip_12_16,x[12],y[16]);
and and785(ip_12_17,x[12],y[17]);
and and786(ip_12_18,x[12],y[18]);
and and787(ip_12_19,x[12],y[19]);
and and788(ip_12_20,x[12],y[20]);
and and789(ip_12_21,x[12],y[21]);
and and790(ip_12_22,x[12],y[22]);
and and791(ip_12_23,x[12],y[23]);
and and792(ip_12_24,x[12],y[24]);
and and793(ip_12_25,x[12],y[25]);
and and794(ip_12_26,x[12],y[26]);
and and795(ip_12_27,x[12],y[27]);
and and796(ip_12_28,x[12],y[28]);
and and797(ip_12_29,x[12],y[29]);
and and798(ip_12_30,x[12],y[30]);
and and799(ip_12_31,x[12],y[31]);
and and800(ip_12_32,x[12],y[32]);
and and801(ip_12_33,x[12],y[33]);
and and802(ip_12_34,x[12],y[34]);
and and803(ip_12_35,x[12],y[35]);
and and804(ip_12_36,x[12],y[36]);
and and805(ip_12_37,x[12],y[37]);
and and806(ip_12_38,x[12],y[38]);
and and807(ip_12_39,x[12],y[39]);
and and808(ip_12_40,x[12],y[40]);
and and809(ip_12_41,x[12],y[41]);
and and810(ip_12_42,x[12],y[42]);
and and811(ip_12_43,x[12],y[43]);
and and812(ip_12_44,x[12],y[44]);
and and813(ip_12_45,x[12],y[45]);
and and814(ip_12_46,x[12],y[46]);
and and815(ip_12_47,x[12],y[47]);
and and816(ip_12_48,x[12],y[48]);
and and817(ip_12_49,x[12],y[49]);
and and818(ip_12_50,x[12],y[50]);
and and819(ip_12_51,x[12],y[51]);
and and820(ip_12_52,x[12],y[52]);
and and821(ip_12_53,x[12],y[53]);
and and822(ip_12_54,x[12],y[54]);
and and823(ip_12_55,x[12],y[55]);
and and824(ip_12_56,x[12],y[56]);
and and825(ip_12_57,x[12],y[57]);
and and826(ip_12_58,x[12],y[58]);
and and827(ip_12_59,x[12],y[59]);
and and828(ip_12_60,x[12],y[60]);
and and829(ip_12_61,x[12],y[61]);
and and830(ip_12_62,x[12],y[62]);
and and831(ip_12_63,x[12],y[63]);
and and832(ip_13_0,x[13],y[0]);
and and833(ip_13_1,x[13],y[1]);
and and834(ip_13_2,x[13],y[2]);
and and835(ip_13_3,x[13],y[3]);
and and836(ip_13_4,x[13],y[4]);
and and837(ip_13_5,x[13],y[5]);
and and838(ip_13_6,x[13],y[6]);
and and839(ip_13_7,x[13],y[7]);
and and840(ip_13_8,x[13],y[8]);
and and841(ip_13_9,x[13],y[9]);
and and842(ip_13_10,x[13],y[10]);
and and843(ip_13_11,x[13],y[11]);
and and844(ip_13_12,x[13],y[12]);
and and845(ip_13_13,x[13],y[13]);
and and846(ip_13_14,x[13],y[14]);
and and847(ip_13_15,x[13],y[15]);
and and848(ip_13_16,x[13],y[16]);
and and849(ip_13_17,x[13],y[17]);
and and850(ip_13_18,x[13],y[18]);
and and851(ip_13_19,x[13],y[19]);
and and852(ip_13_20,x[13],y[20]);
and and853(ip_13_21,x[13],y[21]);
and and854(ip_13_22,x[13],y[22]);
and and855(ip_13_23,x[13],y[23]);
and and856(ip_13_24,x[13],y[24]);
and and857(ip_13_25,x[13],y[25]);
and and858(ip_13_26,x[13],y[26]);
and and859(ip_13_27,x[13],y[27]);
and and860(ip_13_28,x[13],y[28]);
and and861(ip_13_29,x[13],y[29]);
and and862(ip_13_30,x[13],y[30]);
and and863(ip_13_31,x[13],y[31]);
and and864(ip_13_32,x[13],y[32]);
and and865(ip_13_33,x[13],y[33]);
and and866(ip_13_34,x[13],y[34]);
and and867(ip_13_35,x[13],y[35]);
and and868(ip_13_36,x[13],y[36]);
and and869(ip_13_37,x[13],y[37]);
and and870(ip_13_38,x[13],y[38]);
and and871(ip_13_39,x[13],y[39]);
and and872(ip_13_40,x[13],y[40]);
and and873(ip_13_41,x[13],y[41]);
and and874(ip_13_42,x[13],y[42]);
and and875(ip_13_43,x[13],y[43]);
and and876(ip_13_44,x[13],y[44]);
and and877(ip_13_45,x[13],y[45]);
and and878(ip_13_46,x[13],y[46]);
and and879(ip_13_47,x[13],y[47]);
and and880(ip_13_48,x[13],y[48]);
and and881(ip_13_49,x[13],y[49]);
and and882(ip_13_50,x[13],y[50]);
and and883(ip_13_51,x[13],y[51]);
and and884(ip_13_52,x[13],y[52]);
and and885(ip_13_53,x[13],y[53]);
and and886(ip_13_54,x[13],y[54]);
and and887(ip_13_55,x[13],y[55]);
and and888(ip_13_56,x[13],y[56]);
and and889(ip_13_57,x[13],y[57]);
and and890(ip_13_58,x[13],y[58]);
and and891(ip_13_59,x[13],y[59]);
and and892(ip_13_60,x[13],y[60]);
and and893(ip_13_61,x[13],y[61]);
and and894(ip_13_62,x[13],y[62]);
and and895(ip_13_63,x[13],y[63]);
and and896(ip_14_0,x[14],y[0]);
and and897(ip_14_1,x[14],y[1]);
and and898(ip_14_2,x[14],y[2]);
and and899(ip_14_3,x[14],y[3]);
and and900(ip_14_4,x[14],y[4]);
and and901(ip_14_5,x[14],y[5]);
and and902(ip_14_6,x[14],y[6]);
and and903(ip_14_7,x[14],y[7]);
and and904(ip_14_8,x[14],y[8]);
and and905(ip_14_9,x[14],y[9]);
and and906(ip_14_10,x[14],y[10]);
and and907(ip_14_11,x[14],y[11]);
and and908(ip_14_12,x[14],y[12]);
and and909(ip_14_13,x[14],y[13]);
and and910(ip_14_14,x[14],y[14]);
and and911(ip_14_15,x[14],y[15]);
and and912(ip_14_16,x[14],y[16]);
and and913(ip_14_17,x[14],y[17]);
and and914(ip_14_18,x[14],y[18]);
and and915(ip_14_19,x[14],y[19]);
and and916(ip_14_20,x[14],y[20]);
and and917(ip_14_21,x[14],y[21]);
and and918(ip_14_22,x[14],y[22]);
and and919(ip_14_23,x[14],y[23]);
and and920(ip_14_24,x[14],y[24]);
and and921(ip_14_25,x[14],y[25]);
and and922(ip_14_26,x[14],y[26]);
and and923(ip_14_27,x[14],y[27]);
and and924(ip_14_28,x[14],y[28]);
and and925(ip_14_29,x[14],y[29]);
and and926(ip_14_30,x[14],y[30]);
and and927(ip_14_31,x[14],y[31]);
and and928(ip_14_32,x[14],y[32]);
and and929(ip_14_33,x[14],y[33]);
and and930(ip_14_34,x[14],y[34]);
and and931(ip_14_35,x[14],y[35]);
and and932(ip_14_36,x[14],y[36]);
and and933(ip_14_37,x[14],y[37]);
and and934(ip_14_38,x[14],y[38]);
and and935(ip_14_39,x[14],y[39]);
and and936(ip_14_40,x[14],y[40]);
and and937(ip_14_41,x[14],y[41]);
and and938(ip_14_42,x[14],y[42]);
and and939(ip_14_43,x[14],y[43]);
and and940(ip_14_44,x[14],y[44]);
and and941(ip_14_45,x[14],y[45]);
and and942(ip_14_46,x[14],y[46]);
and and943(ip_14_47,x[14],y[47]);
and and944(ip_14_48,x[14],y[48]);
and and945(ip_14_49,x[14],y[49]);
and and946(ip_14_50,x[14],y[50]);
and and947(ip_14_51,x[14],y[51]);
and and948(ip_14_52,x[14],y[52]);
and and949(ip_14_53,x[14],y[53]);
and and950(ip_14_54,x[14],y[54]);
and and951(ip_14_55,x[14],y[55]);
and and952(ip_14_56,x[14],y[56]);
and and953(ip_14_57,x[14],y[57]);
and and954(ip_14_58,x[14],y[58]);
and and955(ip_14_59,x[14],y[59]);
and and956(ip_14_60,x[14],y[60]);
and and957(ip_14_61,x[14],y[61]);
and and958(ip_14_62,x[14],y[62]);
and and959(ip_14_63,x[14],y[63]);
and and960(ip_15_0,x[15],y[0]);
and and961(ip_15_1,x[15],y[1]);
and and962(ip_15_2,x[15],y[2]);
and and963(ip_15_3,x[15],y[3]);
and and964(ip_15_4,x[15],y[4]);
and and965(ip_15_5,x[15],y[5]);
and and966(ip_15_6,x[15],y[6]);
and and967(ip_15_7,x[15],y[7]);
and and968(ip_15_8,x[15],y[8]);
and and969(ip_15_9,x[15],y[9]);
and and970(ip_15_10,x[15],y[10]);
and and971(ip_15_11,x[15],y[11]);
and and972(ip_15_12,x[15],y[12]);
and and973(ip_15_13,x[15],y[13]);
and and974(ip_15_14,x[15],y[14]);
and and975(ip_15_15,x[15],y[15]);
and and976(ip_15_16,x[15],y[16]);
and and977(ip_15_17,x[15],y[17]);
and and978(ip_15_18,x[15],y[18]);
and and979(ip_15_19,x[15],y[19]);
and and980(ip_15_20,x[15],y[20]);
and and981(ip_15_21,x[15],y[21]);
and and982(ip_15_22,x[15],y[22]);
and and983(ip_15_23,x[15],y[23]);
and and984(ip_15_24,x[15],y[24]);
and and985(ip_15_25,x[15],y[25]);
and and986(ip_15_26,x[15],y[26]);
and and987(ip_15_27,x[15],y[27]);
and and988(ip_15_28,x[15],y[28]);
and and989(ip_15_29,x[15],y[29]);
and and990(ip_15_30,x[15],y[30]);
and and991(ip_15_31,x[15],y[31]);
and and992(ip_15_32,x[15],y[32]);
and and993(ip_15_33,x[15],y[33]);
and and994(ip_15_34,x[15],y[34]);
and and995(ip_15_35,x[15],y[35]);
and and996(ip_15_36,x[15],y[36]);
and and997(ip_15_37,x[15],y[37]);
and and998(ip_15_38,x[15],y[38]);
and and999(ip_15_39,x[15],y[39]);
and and1000(ip_15_40,x[15],y[40]);
and and1001(ip_15_41,x[15],y[41]);
and and1002(ip_15_42,x[15],y[42]);
and and1003(ip_15_43,x[15],y[43]);
and and1004(ip_15_44,x[15],y[44]);
and and1005(ip_15_45,x[15],y[45]);
and and1006(ip_15_46,x[15],y[46]);
and and1007(ip_15_47,x[15],y[47]);
and and1008(ip_15_48,x[15],y[48]);
and and1009(ip_15_49,x[15],y[49]);
and and1010(ip_15_50,x[15],y[50]);
and and1011(ip_15_51,x[15],y[51]);
and and1012(ip_15_52,x[15],y[52]);
and and1013(ip_15_53,x[15],y[53]);
and and1014(ip_15_54,x[15],y[54]);
and and1015(ip_15_55,x[15],y[55]);
and and1016(ip_15_56,x[15],y[56]);
and and1017(ip_15_57,x[15],y[57]);
and and1018(ip_15_58,x[15],y[58]);
and and1019(ip_15_59,x[15],y[59]);
and and1020(ip_15_60,x[15],y[60]);
and and1021(ip_15_61,x[15],y[61]);
and and1022(ip_15_62,x[15],y[62]);
and and1023(ip_15_63,x[15],y[63]);
and and1024(ip_16_0,x[16],y[0]);
and and1025(ip_16_1,x[16],y[1]);
and and1026(ip_16_2,x[16],y[2]);
and and1027(ip_16_3,x[16],y[3]);
and and1028(ip_16_4,x[16],y[4]);
and and1029(ip_16_5,x[16],y[5]);
and and1030(ip_16_6,x[16],y[6]);
and and1031(ip_16_7,x[16],y[7]);
and and1032(ip_16_8,x[16],y[8]);
and and1033(ip_16_9,x[16],y[9]);
and and1034(ip_16_10,x[16],y[10]);
and and1035(ip_16_11,x[16],y[11]);
and and1036(ip_16_12,x[16],y[12]);
and and1037(ip_16_13,x[16],y[13]);
and and1038(ip_16_14,x[16],y[14]);
and and1039(ip_16_15,x[16],y[15]);
and and1040(ip_16_16,x[16],y[16]);
and and1041(ip_16_17,x[16],y[17]);
and and1042(ip_16_18,x[16],y[18]);
and and1043(ip_16_19,x[16],y[19]);
and and1044(ip_16_20,x[16],y[20]);
and and1045(ip_16_21,x[16],y[21]);
and and1046(ip_16_22,x[16],y[22]);
and and1047(ip_16_23,x[16],y[23]);
and and1048(ip_16_24,x[16],y[24]);
and and1049(ip_16_25,x[16],y[25]);
and and1050(ip_16_26,x[16],y[26]);
and and1051(ip_16_27,x[16],y[27]);
and and1052(ip_16_28,x[16],y[28]);
and and1053(ip_16_29,x[16],y[29]);
and and1054(ip_16_30,x[16],y[30]);
and and1055(ip_16_31,x[16],y[31]);
and and1056(ip_16_32,x[16],y[32]);
and and1057(ip_16_33,x[16],y[33]);
and and1058(ip_16_34,x[16],y[34]);
and and1059(ip_16_35,x[16],y[35]);
and and1060(ip_16_36,x[16],y[36]);
and and1061(ip_16_37,x[16],y[37]);
and and1062(ip_16_38,x[16],y[38]);
and and1063(ip_16_39,x[16],y[39]);
and and1064(ip_16_40,x[16],y[40]);
and and1065(ip_16_41,x[16],y[41]);
and and1066(ip_16_42,x[16],y[42]);
and and1067(ip_16_43,x[16],y[43]);
and and1068(ip_16_44,x[16],y[44]);
and and1069(ip_16_45,x[16],y[45]);
and and1070(ip_16_46,x[16],y[46]);
and and1071(ip_16_47,x[16],y[47]);
and and1072(ip_16_48,x[16],y[48]);
and and1073(ip_16_49,x[16],y[49]);
and and1074(ip_16_50,x[16],y[50]);
and and1075(ip_16_51,x[16],y[51]);
and and1076(ip_16_52,x[16],y[52]);
and and1077(ip_16_53,x[16],y[53]);
and and1078(ip_16_54,x[16],y[54]);
and and1079(ip_16_55,x[16],y[55]);
and and1080(ip_16_56,x[16],y[56]);
and and1081(ip_16_57,x[16],y[57]);
and and1082(ip_16_58,x[16],y[58]);
and and1083(ip_16_59,x[16],y[59]);
and and1084(ip_16_60,x[16],y[60]);
and and1085(ip_16_61,x[16],y[61]);
and and1086(ip_16_62,x[16],y[62]);
and and1087(ip_16_63,x[16],y[63]);
and and1088(ip_17_0,x[17],y[0]);
and and1089(ip_17_1,x[17],y[1]);
and and1090(ip_17_2,x[17],y[2]);
and and1091(ip_17_3,x[17],y[3]);
and and1092(ip_17_4,x[17],y[4]);
and and1093(ip_17_5,x[17],y[5]);
and and1094(ip_17_6,x[17],y[6]);
and and1095(ip_17_7,x[17],y[7]);
and and1096(ip_17_8,x[17],y[8]);
and and1097(ip_17_9,x[17],y[9]);
and and1098(ip_17_10,x[17],y[10]);
and and1099(ip_17_11,x[17],y[11]);
and and1100(ip_17_12,x[17],y[12]);
and and1101(ip_17_13,x[17],y[13]);
and and1102(ip_17_14,x[17],y[14]);
and and1103(ip_17_15,x[17],y[15]);
and and1104(ip_17_16,x[17],y[16]);
and and1105(ip_17_17,x[17],y[17]);
and and1106(ip_17_18,x[17],y[18]);
and and1107(ip_17_19,x[17],y[19]);
and and1108(ip_17_20,x[17],y[20]);
and and1109(ip_17_21,x[17],y[21]);
and and1110(ip_17_22,x[17],y[22]);
and and1111(ip_17_23,x[17],y[23]);
and and1112(ip_17_24,x[17],y[24]);
and and1113(ip_17_25,x[17],y[25]);
and and1114(ip_17_26,x[17],y[26]);
and and1115(ip_17_27,x[17],y[27]);
and and1116(ip_17_28,x[17],y[28]);
and and1117(ip_17_29,x[17],y[29]);
and and1118(ip_17_30,x[17],y[30]);
and and1119(ip_17_31,x[17],y[31]);
and and1120(ip_17_32,x[17],y[32]);
and and1121(ip_17_33,x[17],y[33]);
and and1122(ip_17_34,x[17],y[34]);
and and1123(ip_17_35,x[17],y[35]);
and and1124(ip_17_36,x[17],y[36]);
and and1125(ip_17_37,x[17],y[37]);
and and1126(ip_17_38,x[17],y[38]);
and and1127(ip_17_39,x[17],y[39]);
and and1128(ip_17_40,x[17],y[40]);
and and1129(ip_17_41,x[17],y[41]);
and and1130(ip_17_42,x[17],y[42]);
and and1131(ip_17_43,x[17],y[43]);
and and1132(ip_17_44,x[17],y[44]);
and and1133(ip_17_45,x[17],y[45]);
and and1134(ip_17_46,x[17],y[46]);
and and1135(ip_17_47,x[17],y[47]);
and and1136(ip_17_48,x[17],y[48]);
and and1137(ip_17_49,x[17],y[49]);
and and1138(ip_17_50,x[17],y[50]);
and and1139(ip_17_51,x[17],y[51]);
and and1140(ip_17_52,x[17],y[52]);
and and1141(ip_17_53,x[17],y[53]);
and and1142(ip_17_54,x[17],y[54]);
and and1143(ip_17_55,x[17],y[55]);
and and1144(ip_17_56,x[17],y[56]);
and and1145(ip_17_57,x[17],y[57]);
and and1146(ip_17_58,x[17],y[58]);
and and1147(ip_17_59,x[17],y[59]);
and and1148(ip_17_60,x[17],y[60]);
and and1149(ip_17_61,x[17],y[61]);
and and1150(ip_17_62,x[17],y[62]);
and and1151(ip_17_63,x[17],y[63]);
and and1152(ip_18_0,x[18],y[0]);
and and1153(ip_18_1,x[18],y[1]);
and and1154(ip_18_2,x[18],y[2]);
and and1155(ip_18_3,x[18],y[3]);
and and1156(ip_18_4,x[18],y[4]);
and and1157(ip_18_5,x[18],y[5]);
and and1158(ip_18_6,x[18],y[6]);
and and1159(ip_18_7,x[18],y[7]);
and and1160(ip_18_8,x[18],y[8]);
and and1161(ip_18_9,x[18],y[9]);
and and1162(ip_18_10,x[18],y[10]);
and and1163(ip_18_11,x[18],y[11]);
and and1164(ip_18_12,x[18],y[12]);
and and1165(ip_18_13,x[18],y[13]);
and and1166(ip_18_14,x[18],y[14]);
and and1167(ip_18_15,x[18],y[15]);
and and1168(ip_18_16,x[18],y[16]);
and and1169(ip_18_17,x[18],y[17]);
and and1170(ip_18_18,x[18],y[18]);
and and1171(ip_18_19,x[18],y[19]);
and and1172(ip_18_20,x[18],y[20]);
and and1173(ip_18_21,x[18],y[21]);
and and1174(ip_18_22,x[18],y[22]);
and and1175(ip_18_23,x[18],y[23]);
and and1176(ip_18_24,x[18],y[24]);
and and1177(ip_18_25,x[18],y[25]);
and and1178(ip_18_26,x[18],y[26]);
and and1179(ip_18_27,x[18],y[27]);
and and1180(ip_18_28,x[18],y[28]);
and and1181(ip_18_29,x[18],y[29]);
and and1182(ip_18_30,x[18],y[30]);
and and1183(ip_18_31,x[18],y[31]);
and and1184(ip_18_32,x[18],y[32]);
and and1185(ip_18_33,x[18],y[33]);
and and1186(ip_18_34,x[18],y[34]);
and and1187(ip_18_35,x[18],y[35]);
and and1188(ip_18_36,x[18],y[36]);
and and1189(ip_18_37,x[18],y[37]);
and and1190(ip_18_38,x[18],y[38]);
and and1191(ip_18_39,x[18],y[39]);
and and1192(ip_18_40,x[18],y[40]);
and and1193(ip_18_41,x[18],y[41]);
and and1194(ip_18_42,x[18],y[42]);
and and1195(ip_18_43,x[18],y[43]);
and and1196(ip_18_44,x[18],y[44]);
and and1197(ip_18_45,x[18],y[45]);
and and1198(ip_18_46,x[18],y[46]);
and and1199(ip_18_47,x[18],y[47]);
and and1200(ip_18_48,x[18],y[48]);
and and1201(ip_18_49,x[18],y[49]);
and and1202(ip_18_50,x[18],y[50]);
and and1203(ip_18_51,x[18],y[51]);
and and1204(ip_18_52,x[18],y[52]);
and and1205(ip_18_53,x[18],y[53]);
and and1206(ip_18_54,x[18],y[54]);
and and1207(ip_18_55,x[18],y[55]);
and and1208(ip_18_56,x[18],y[56]);
and and1209(ip_18_57,x[18],y[57]);
and and1210(ip_18_58,x[18],y[58]);
and and1211(ip_18_59,x[18],y[59]);
and and1212(ip_18_60,x[18],y[60]);
and and1213(ip_18_61,x[18],y[61]);
and and1214(ip_18_62,x[18],y[62]);
and and1215(ip_18_63,x[18],y[63]);
and and1216(ip_19_0,x[19],y[0]);
and and1217(ip_19_1,x[19],y[1]);
and and1218(ip_19_2,x[19],y[2]);
and and1219(ip_19_3,x[19],y[3]);
and and1220(ip_19_4,x[19],y[4]);
and and1221(ip_19_5,x[19],y[5]);
and and1222(ip_19_6,x[19],y[6]);
and and1223(ip_19_7,x[19],y[7]);
and and1224(ip_19_8,x[19],y[8]);
and and1225(ip_19_9,x[19],y[9]);
and and1226(ip_19_10,x[19],y[10]);
and and1227(ip_19_11,x[19],y[11]);
and and1228(ip_19_12,x[19],y[12]);
and and1229(ip_19_13,x[19],y[13]);
and and1230(ip_19_14,x[19],y[14]);
and and1231(ip_19_15,x[19],y[15]);
and and1232(ip_19_16,x[19],y[16]);
and and1233(ip_19_17,x[19],y[17]);
and and1234(ip_19_18,x[19],y[18]);
and and1235(ip_19_19,x[19],y[19]);
and and1236(ip_19_20,x[19],y[20]);
and and1237(ip_19_21,x[19],y[21]);
and and1238(ip_19_22,x[19],y[22]);
and and1239(ip_19_23,x[19],y[23]);
and and1240(ip_19_24,x[19],y[24]);
and and1241(ip_19_25,x[19],y[25]);
and and1242(ip_19_26,x[19],y[26]);
and and1243(ip_19_27,x[19],y[27]);
and and1244(ip_19_28,x[19],y[28]);
and and1245(ip_19_29,x[19],y[29]);
and and1246(ip_19_30,x[19],y[30]);
and and1247(ip_19_31,x[19],y[31]);
and and1248(ip_19_32,x[19],y[32]);
and and1249(ip_19_33,x[19],y[33]);
and and1250(ip_19_34,x[19],y[34]);
and and1251(ip_19_35,x[19],y[35]);
and and1252(ip_19_36,x[19],y[36]);
and and1253(ip_19_37,x[19],y[37]);
and and1254(ip_19_38,x[19],y[38]);
and and1255(ip_19_39,x[19],y[39]);
and and1256(ip_19_40,x[19],y[40]);
and and1257(ip_19_41,x[19],y[41]);
and and1258(ip_19_42,x[19],y[42]);
and and1259(ip_19_43,x[19],y[43]);
and and1260(ip_19_44,x[19],y[44]);
and and1261(ip_19_45,x[19],y[45]);
and and1262(ip_19_46,x[19],y[46]);
and and1263(ip_19_47,x[19],y[47]);
and and1264(ip_19_48,x[19],y[48]);
and and1265(ip_19_49,x[19],y[49]);
and and1266(ip_19_50,x[19],y[50]);
and and1267(ip_19_51,x[19],y[51]);
and and1268(ip_19_52,x[19],y[52]);
and and1269(ip_19_53,x[19],y[53]);
and and1270(ip_19_54,x[19],y[54]);
and and1271(ip_19_55,x[19],y[55]);
and and1272(ip_19_56,x[19],y[56]);
and and1273(ip_19_57,x[19],y[57]);
and and1274(ip_19_58,x[19],y[58]);
and and1275(ip_19_59,x[19],y[59]);
and and1276(ip_19_60,x[19],y[60]);
and and1277(ip_19_61,x[19],y[61]);
and and1278(ip_19_62,x[19],y[62]);
and and1279(ip_19_63,x[19],y[63]);
and and1280(ip_20_0,x[20],y[0]);
and and1281(ip_20_1,x[20],y[1]);
and and1282(ip_20_2,x[20],y[2]);
and and1283(ip_20_3,x[20],y[3]);
and and1284(ip_20_4,x[20],y[4]);
and and1285(ip_20_5,x[20],y[5]);
and and1286(ip_20_6,x[20],y[6]);
and and1287(ip_20_7,x[20],y[7]);
and and1288(ip_20_8,x[20],y[8]);
and and1289(ip_20_9,x[20],y[9]);
and and1290(ip_20_10,x[20],y[10]);
and and1291(ip_20_11,x[20],y[11]);
and and1292(ip_20_12,x[20],y[12]);
and and1293(ip_20_13,x[20],y[13]);
and and1294(ip_20_14,x[20],y[14]);
and and1295(ip_20_15,x[20],y[15]);
and and1296(ip_20_16,x[20],y[16]);
and and1297(ip_20_17,x[20],y[17]);
and and1298(ip_20_18,x[20],y[18]);
and and1299(ip_20_19,x[20],y[19]);
and and1300(ip_20_20,x[20],y[20]);
and and1301(ip_20_21,x[20],y[21]);
and and1302(ip_20_22,x[20],y[22]);
and and1303(ip_20_23,x[20],y[23]);
and and1304(ip_20_24,x[20],y[24]);
and and1305(ip_20_25,x[20],y[25]);
and and1306(ip_20_26,x[20],y[26]);
and and1307(ip_20_27,x[20],y[27]);
and and1308(ip_20_28,x[20],y[28]);
and and1309(ip_20_29,x[20],y[29]);
and and1310(ip_20_30,x[20],y[30]);
and and1311(ip_20_31,x[20],y[31]);
and and1312(ip_20_32,x[20],y[32]);
and and1313(ip_20_33,x[20],y[33]);
and and1314(ip_20_34,x[20],y[34]);
and and1315(ip_20_35,x[20],y[35]);
and and1316(ip_20_36,x[20],y[36]);
and and1317(ip_20_37,x[20],y[37]);
and and1318(ip_20_38,x[20],y[38]);
and and1319(ip_20_39,x[20],y[39]);
and and1320(ip_20_40,x[20],y[40]);
and and1321(ip_20_41,x[20],y[41]);
and and1322(ip_20_42,x[20],y[42]);
and and1323(ip_20_43,x[20],y[43]);
and and1324(ip_20_44,x[20],y[44]);
and and1325(ip_20_45,x[20],y[45]);
and and1326(ip_20_46,x[20],y[46]);
and and1327(ip_20_47,x[20],y[47]);
and and1328(ip_20_48,x[20],y[48]);
and and1329(ip_20_49,x[20],y[49]);
and and1330(ip_20_50,x[20],y[50]);
and and1331(ip_20_51,x[20],y[51]);
and and1332(ip_20_52,x[20],y[52]);
and and1333(ip_20_53,x[20],y[53]);
and and1334(ip_20_54,x[20],y[54]);
and and1335(ip_20_55,x[20],y[55]);
and and1336(ip_20_56,x[20],y[56]);
and and1337(ip_20_57,x[20],y[57]);
and and1338(ip_20_58,x[20],y[58]);
and and1339(ip_20_59,x[20],y[59]);
and and1340(ip_20_60,x[20],y[60]);
and and1341(ip_20_61,x[20],y[61]);
and and1342(ip_20_62,x[20],y[62]);
and and1343(ip_20_63,x[20],y[63]);
and and1344(ip_21_0,x[21],y[0]);
and and1345(ip_21_1,x[21],y[1]);
and and1346(ip_21_2,x[21],y[2]);
and and1347(ip_21_3,x[21],y[3]);
and and1348(ip_21_4,x[21],y[4]);
and and1349(ip_21_5,x[21],y[5]);
and and1350(ip_21_6,x[21],y[6]);
and and1351(ip_21_7,x[21],y[7]);
and and1352(ip_21_8,x[21],y[8]);
and and1353(ip_21_9,x[21],y[9]);
and and1354(ip_21_10,x[21],y[10]);
and and1355(ip_21_11,x[21],y[11]);
and and1356(ip_21_12,x[21],y[12]);
and and1357(ip_21_13,x[21],y[13]);
and and1358(ip_21_14,x[21],y[14]);
and and1359(ip_21_15,x[21],y[15]);
and and1360(ip_21_16,x[21],y[16]);
and and1361(ip_21_17,x[21],y[17]);
and and1362(ip_21_18,x[21],y[18]);
and and1363(ip_21_19,x[21],y[19]);
and and1364(ip_21_20,x[21],y[20]);
and and1365(ip_21_21,x[21],y[21]);
and and1366(ip_21_22,x[21],y[22]);
and and1367(ip_21_23,x[21],y[23]);
and and1368(ip_21_24,x[21],y[24]);
and and1369(ip_21_25,x[21],y[25]);
and and1370(ip_21_26,x[21],y[26]);
and and1371(ip_21_27,x[21],y[27]);
and and1372(ip_21_28,x[21],y[28]);
and and1373(ip_21_29,x[21],y[29]);
and and1374(ip_21_30,x[21],y[30]);
and and1375(ip_21_31,x[21],y[31]);
and and1376(ip_21_32,x[21],y[32]);
and and1377(ip_21_33,x[21],y[33]);
and and1378(ip_21_34,x[21],y[34]);
and and1379(ip_21_35,x[21],y[35]);
and and1380(ip_21_36,x[21],y[36]);
and and1381(ip_21_37,x[21],y[37]);
and and1382(ip_21_38,x[21],y[38]);
and and1383(ip_21_39,x[21],y[39]);
and and1384(ip_21_40,x[21],y[40]);
and and1385(ip_21_41,x[21],y[41]);
and and1386(ip_21_42,x[21],y[42]);
and and1387(ip_21_43,x[21],y[43]);
and and1388(ip_21_44,x[21],y[44]);
and and1389(ip_21_45,x[21],y[45]);
and and1390(ip_21_46,x[21],y[46]);
and and1391(ip_21_47,x[21],y[47]);
and and1392(ip_21_48,x[21],y[48]);
and and1393(ip_21_49,x[21],y[49]);
and and1394(ip_21_50,x[21],y[50]);
and and1395(ip_21_51,x[21],y[51]);
and and1396(ip_21_52,x[21],y[52]);
and and1397(ip_21_53,x[21],y[53]);
and and1398(ip_21_54,x[21],y[54]);
and and1399(ip_21_55,x[21],y[55]);
and and1400(ip_21_56,x[21],y[56]);
and and1401(ip_21_57,x[21],y[57]);
and and1402(ip_21_58,x[21],y[58]);
and and1403(ip_21_59,x[21],y[59]);
and and1404(ip_21_60,x[21],y[60]);
and and1405(ip_21_61,x[21],y[61]);
and and1406(ip_21_62,x[21],y[62]);
and and1407(ip_21_63,x[21],y[63]);
and and1408(ip_22_0,x[22],y[0]);
and and1409(ip_22_1,x[22],y[1]);
and and1410(ip_22_2,x[22],y[2]);
and and1411(ip_22_3,x[22],y[3]);
and and1412(ip_22_4,x[22],y[4]);
and and1413(ip_22_5,x[22],y[5]);
and and1414(ip_22_6,x[22],y[6]);
and and1415(ip_22_7,x[22],y[7]);
and and1416(ip_22_8,x[22],y[8]);
and and1417(ip_22_9,x[22],y[9]);
and and1418(ip_22_10,x[22],y[10]);
and and1419(ip_22_11,x[22],y[11]);
and and1420(ip_22_12,x[22],y[12]);
and and1421(ip_22_13,x[22],y[13]);
and and1422(ip_22_14,x[22],y[14]);
and and1423(ip_22_15,x[22],y[15]);
and and1424(ip_22_16,x[22],y[16]);
and and1425(ip_22_17,x[22],y[17]);
and and1426(ip_22_18,x[22],y[18]);
and and1427(ip_22_19,x[22],y[19]);
and and1428(ip_22_20,x[22],y[20]);
and and1429(ip_22_21,x[22],y[21]);
and and1430(ip_22_22,x[22],y[22]);
and and1431(ip_22_23,x[22],y[23]);
and and1432(ip_22_24,x[22],y[24]);
and and1433(ip_22_25,x[22],y[25]);
and and1434(ip_22_26,x[22],y[26]);
and and1435(ip_22_27,x[22],y[27]);
and and1436(ip_22_28,x[22],y[28]);
and and1437(ip_22_29,x[22],y[29]);
and and1438(ip_22_30,x[22],y[30]);
and and1439(ip_22_31,x[22],y[31]);
and and1440(ip_22_32,x[22],y[32]);
and and1441(ip_22_33,x[22],y[33]);
and and1442(ip_22_34,x[22],y[34]);
and and1443(ip_22_35,x[22],y[35]);
and and1444(ip_22_36,x[22],y[36]);
and and1445(ip_22_37,x[22],y[37]);
and and1446(ip_22_38,x[22],y[38]);
and and1447(ip_22_39,x[22],y[39]);
and and1448(ip_22_40,x[22],y[40]);
and and1449(ip_22_41,x[22],y[41]);
and and1450(ip_22_42,x[22],y[42]);
and and1451(ip_22_43,x[22],y[43]);
and and1452(ip_22_44,x[22],y[44]);
and and1453(ip_22_45,x[22],y[45]);
and and1454(ip_22_46,x[22],y[46]);
and and1455(ip_22_47,x[22],y[47]);
and and1456(ip_22_48,x[22],y[48]);
and and1457(ip_22_49,x[22],y[49]);
and and1458(ip_22_50,x[22],y[50]);
and and1459(ip_22_51,x[22],y[51]);
and and1460(ip_22_52,x[22],y[52]);
and and1461(ip_22_53,x[22],y[53]);
and and1462(ip_22_54,x[22],y[54]);
and and1463(ip_22_55,x[22],y[55]);
and and1464(ip_22_56,x[22],y[56]);
and and1465(ip_22_57,x[22],y[57]);
and and1466(ip_22_58,x[22],y[58]);
and and1467(ip_22_59,x[22],y[59]);
and and1468(ip_22_60,x[22],y[60]);
and and1469(ip_22_61,x[22],y[61]);
and and1470(ip_22_62,x[22],y[62]);
and and1471(ip_22_63,x[22],y[63]);
and and1472(ip_23_0,x[23],y[0]);
and and1473(ip_23_1,x[23],y[1]);
and and1474(ip_23_2,x[23],y[2]);
and and1475(ip_23_3,x[23],y[3]);
and and1476(ip_23_4,x[23],y[4]);
and and1477(ip_23_5,x[23],y[5]);
and and1478(ip_23_6,x[23],y[6]);
and and1479(ip_23_7,x[23],y[7]);
and and1480(ip_23_8,x[23],y[8]);
and and1481(ip_23_9,x[23],y[9]);
and and1482(ip_23_10,x[23],y[10]);
and and1483(ip_23_11,x[23],y[11]);
and and1484(ip_23_12,x[23],y[12]);
and and1485(ip_23_13,x[23],y[13]);
and and1486(ip_23_14,x[23],y[14]);
and and1487(ip_23_15,x[23],y[15]);
and and1488(ip_23_16,x[23],y[16]);
and and1489(ip_23_17,x[23],y[17]);
and and1490(ip_23_18,x[23],y[18]);
and and1491(ip_23_19,x[23],y[19]);
and and1492(ip_23_20,x[23],y[20]);
and and1493(ip_23_21,x[23],y[21]);
and and1494(ip_23_22,x[23],y[22]);
and and1495(ip_23_23,x[23],y[23]);
and and1496(ip_23_24,x[23],y[24]);
and and1497(ip_23_25,x[23],y[25]);
and and1498(ip_23_26,x[23],y[26]);
and and1499(ip_23_27,x[23],y[27]);
and and1500(ip_23_28,x[23],y[28]);
and and1501(ip_23_29,x[23],y[29]);
and and1502(ip_23_30,x[23],y[30]);
and and1503(ip_23_31,x[23],y[31]);
and and1504(ip_23_32,x[23],y[32]);
and and1505(ip_23_33,x[23],y[33]);
and and1506(ip_23_34,x[23],y[34]);
and and1507(ip_23_35,x[23],y[35]);
and and1508(ip_23_36,x[23],y[36]);
and and1509(ip_23_37,x[23],y[37]);
and and1510(ip_23_38,x[23],y[38]);
and and1511(ip_23_39,x[23],y[39]);
and and1512(ip_23_40,x[23],y[40]);
and and1513(ip_23_41,x[23],y[41]);
and and1514(ip_23_42,x[23],y[42]);
and and1515(ip_23_43,x[23],y[43]);
and and1516(ip_23_44,x[23],y[44]);
and and1517(ip_23_45,x[23],y[45]);
and and1518(ip_23_46,x[23],y[46]);
and and1519(ip_23_47,x[23],y[47]);
and and1520(ip_23_48,x[23],y[48]);
and and1521(ip_23_49,x[23],y[49]);
and and1522(ip_23_50,x[23],y[50]);
and and1523(ip_23_51,x[23],y[51]);
and and1524(ip_23_52,x[23],y[52]);
and and1525(ip_23_53,x[23],y[53]);
and and1526(ip_23_54,x[23],y[54]);
and and1527(ip_23_55,x[23],y[55]);
and and1528(ip_23_56,x[23],y[56]);
and and1529(ip_23_57,x[23],y[57]);
and and1530(ip_23_58,x[23],y[58]);
and and1531(ip_23_59,x[23],y[59]);
and and1532(ip_23_60,x[23],y[60]);
and and1533(ip_23_61,x[23],y[61]);
and and1534(ip_23_62,x[23],y[62]);
and and1535(ip_23_63,x[23],y[63]);
and and1536(ip_24_0,x[24],y[0]);
and and1537(ip_24_1,x[24],y[1]);
and and1538(ip_24_2,x[24],y[2]);
and and1539(ip_24_3,x[24],y[3]);
and and1540(ip_24_4,x[24],y[4]);
and and1541(ip_24_5,x[24],y[5]);
and and1542(ip_24_6,x[24],y[6]);
and and1543(ip_24_7,x[24],y[7]);
and and1544(ip_24_8,x[24],y[8]);
and and1545(ip_24_9,x[24],y[9]);
and and1546(ip_24_10,x[24],y[10]);
and and1547(ip_24_11,x[24],y[11]);
and and1548(ip_24_12,x[24],y[12]);
and and1549(ip_24_13,x[24],y[13]);
and and1550(ip_24_14,x[24],y[14]);
and and1551(ip_24_15,x[24],y[15]);
and and1552(ip_24_16,x[24],y[16]);
and and1553(ip_24_17,x[24],y[17]);
and and1554(ip_24_18,x[24],y[18]);
and and1555(ip_24_19,x[24],y[19]);
and and1556(ip_24_20,x[24],y[20]);
and and1557(ip_24_21,x[24],y[21]);
and and1558(ip_24_22,x[24],y[22]);
and and1559(ip_24_23,x[24],y[23]);
and and1560(ip_24_24,x[24],y[24]);
and and1561(ip_24_25,x[24],y[25]);
and and1562(ip_24_26,x[24],y[26]);
and and1563(ip_24_27,x[24],y[27]);
and and1564(ip_24_28,x[24],y[28]);
and and1565(ip_24_29,x[24],y[29]);
and and1566(ip_24_30,x[24],y[30]);
and and1567(ip_24_31,x[24],y[31]);
and and1568(ip_24_32,x[24],y[32]);
and and1569(ip_24_33,x[24],y[33]);
and and1570(ip_24_34,x[24],y[34]);
and and1571(ip_24_35,x[24],y[35]);
and and1572(ip_24_36,x[24],y[36]);
and and1573(ip_24_37,x[24],y[37]);
and and1574(ip_24_38,x[24],y[38]);
and and1575(ip_24_39,x[24],y[39]);
and and1576(ip_24_40,x[24],y[40]);
and and1577(ip_24_41,x[24],y[41]);
and and1578(ip_24_42,x[24],y[42]);
and and1579(ip_24_43,x[24],y[43]);
and and1580(ip_24_44,x[24],y[44]);
and and1581(ip_24_45,x[24],y[45]);
and and1582(ip_24_46,x[24],y[46]);
and and1583(ip_24_47,x[24],y[47]);
and and1584(ip_24_48,x[24],y[48]);
and and1585(ip_24_49,x[24],y[49]);
and and1586(ip_24_50,x[24],y[50]);
and and1587(ip_24_51,x[24],y[51]);
and and1588(ip_24_52,x[24],y[52]);
and and1589(ip_24_53,x[24],y[53]);
and and1590(ip_24_54,x[24],y[54]);
and and1591(ip_24_55,x[24],y[55]);
and and1592(ip_24_56,x[24],y[56]);
and and1593(ip_24_57,x[24],y[57]);
and and1594(ip_24_58,x[24],y[58]);
and and1595(ip_24_59,x[24],y[59]);
and and1596(ip_24_60,x[24],y[60]);
and and1597(ip_24_61,x[24],y[61]);
and and1598(ip_24_62,x[24],y[62]);
and and1599(ip_24_63,x[24],y[63]);
and and1600(ip_25_0,x[25],y[0]);
and and1601(ip_25_1,x[25],y[1]);
and and1602(ip_25_2,x[25],y[2]);
and and1603(ip_25_3,x[25],y[3]);
and and1604(ip_25_4,x[25],y[4]);
and and1605(ip_25_5,x[25],y[5]);
and and1606(ip_25_6,x[25],y[6]);
and and1607(ip_25_7,x[25],y[7]);
and and1608(ip_25_8,x[25],y[8]);
and and1609(ip_25_9,x[25],y[9]);
and and1610(ip_25_10,x[25],y[10]);
and and1611(ip_25_11,x[25],y[11]);
and and1612(ip_25_12,x[25],y[12]);
and and1613(ip_25_13,x[25],y[13]);
and and1614(ip_25_14,x[25],y[14]);
and and1615(ip_25_15,x[25],y[15]);
and and1616(ip_25_16,x[25],y[16]);
and and1617(ip_25_17,x[25],y[17]);
and and1618(ip_25_18,x[25],y[18]);
and and1619(ip_25_19,x[25],y[19]);
and and1620(ip_25_20,x[25],y[20]);
and and1621(ip_25_21,x[25],y[21]);
and and1622(ip_25_22,x[25],y[22]);
and and1623(ip_25_23,x[25],y[23]);
and and1624(ip_25_24,x[25],y[24]);
and and1625(ip_25_25,x[25],y[25]);
and and1626(ip_25_26,x[25],y[26]);
and and1627(ip_25_27,x[25],y[27]);
and and1628(ip_25_28,x[25],y[28]);
and and1629(ip_25_29,x[25],y[29]);
and and1630(ip_25_30,x[25],y[30]);
and and1631(ip_25_31,x[25],y[31]);
and and1632(ip_25_32,x[25],y[32]);
and and1633(ip_25_33,x[25],y[33]);
and and1634(ip_25_34,x[25],y[34]);
and and1635(ip_25_35,x[25],y[35]);
and and1636(ip_25_36,x[25],y[36]);
and and1637(ip_25_37,x[25],y[37]);
and and1638(ip_25_38,x[25],y[38]);
and and1639(ip_25_39,x[25],y[39]);
and and1640(ip_25_40,x[25],y[40]);
and and1641(ip_25_41,x[25],y[41]);
and and1642(ip_25_42,x[25],y[42]);
and and1643(ip_25_43,x[25],y[43]);
and and1644(ip_25_44,x[25],y[44]);
and and1645(ip_25_45,x[25],y[45]);
and and1646(ip_25_46,x[25],y[46]);
and and1647(ip_25_47,x[25],y[47]);
and and1648(ip_25_48,x[25],y[48]);
and and1649(ip_25_49,x[25],y[49]);
and and1650(ip_25_50,x[25],y[50]);
and and1651(ip_25_51,x[25],y[51]);
and and1652(ip_25_52,x[25],y[52]);
and and1653(ip_25_53,x[25],y[53]);
and and1654(ip_25_54,x[25],y[54]);
and and1655(ip_25_55,x[25],y[55]);
and and1656(ip_25_56,x[25],y[56]);
and and1657(ip_25_57,x[25],y[57]);
and and1658(ip_25_58,x[25],y[58]);
and and1659(ip_25_59,x[25],y[59]);
and and1660(ip_25_60,x[25],y[60]);
and and1661(ip_25_61,x[25],y[61]);
and and1662(ip_25_62,x[25],y[62]);
and and1663(ip_25_63,x[25],y[63]);
and and1664(ip_26_0,x[26],y[0]);
and and1665(ip_26_1,x[26],y[1]);
and and1666(ip_26_2,x[26],y[2]);
and and1667(ip_26_3,x[26],y[3]);
and and1668(ip_26_4,x[26],y[4]);
and and1669(ip_26_5,x[26],y[5]);
and and1670(ip_26_6,x[26],y[6]);
and and1671(ip_26_7,x[26],y[7]);
and and1672(ip_26_8,x[26],y[8]);
and and1673(ip_26_9,x[26],y[9]);
and and1674(ip_26_10,x[26],y[10]);
and and1675(ip_26_11,x[26],y[11]);
and and1676(ip_26_12,x[26],y[12]);
and and1677(ip_26_13,x[26],y[13]);
and and1678(ip_26_14,x[26],y[14]);
and and1679(ip_26_15,x[26],y[15]);
and and1680(ip_26_16,x[26],y[16]);
and and1681(ip_26_17,x[26],y[17]);
and and1682(ip_26_18,x[26],y[18]);
and and1683(ip_26_19,x[26],y[19]);
and and1684(ip_26_20,x[26],y[20]);
and and1685(ip_26_21,x[26],y[21]);
and and1686(ip_26_22,x[26],y[22]);
and and1687(ip_26_23,x[26],y[23]);
and and1688(ip_26_24,x[26],y[24]);
and and1689(ip_26_25,x[26],y[25]);
and and1690(ip_26_26,x[26],y[26]);
and and1691(ip_26_27,x[26],y[27]);
and and1692(ip_26_28,x[26],y[28]);
and and1693(ip_26_29,x[26],y[29]);
and and1694(ip_26_30,x[26],y[30]);
and and1695(ip_26_31,x[26],y[31]);
and and1696(ip_26_32,x[26],y[32]);
and and1697(ip_26_33,x[26],y[33]);
and and1698(ip_26_34,x[26],y[34]);
and and1699(ip_26_35,x[26],y[35]);
and and1700(ip_26_36,x[26],y[36]);
and and1701(ip_26_37,x[26],y[37]);
and and1702(ip_26_38,x[26],y[38]);
and and1703(ip_26_39,x[26],y[39]);
and and1704(ip_26_40,x[26],y[40]);
and and1705(ip_26_41,x[26],y[41]);
and and1706(ip_26_42,x[26],y[42]);
and and1707(ip_26_43,x[26],y[43]);
and and1708(ip_26_44,x[26],y[44]);
and and1709(ip_26_45,x[26],y[45]);
and and1710(ip_26_46,x[26],y[46]);
and and1711(ip_26_47,x[26],y[47]);
and and1712(ip_26_48,x[26],y[48]);
and and1713(ip_26_49,x[26],y[49]);
and and1714(ip_26_50,x[26],y[50]);
and and1715(ip_26_51,x[26],y[51]);
and and1716(ip_26_52,x[26],y[52]);
and and1717(ip_26_53,x[26],y[53]);
and and1718(ip_26_54,x[26],y[54]);
and and1719(ip_26_55,x[26],y[55]);
and and1720(ip_26_56,x[26],y[56]);
and and1721(ip_26_57,x[26],y[57]);
and and1722(ip_26_58,x[26],y[58]);
and and1723(ip_26_59,x[26],y[59]);
and and1724(ip_26_60,x[26],y[60]);
and and1725(ip_26_61,x[26],y[61]);
and and1726(ip_26_62,x[26],y[62]);
and and1727(ip_26_63,x[26],y[63]);
and and1728(ip_27_0,x[27],y[0]);
and and1729(ip_27_1,x[27],y[1]);
and and1730(ip_27_2,x[27],y[2]);
and and1731(ip_27_3,x[27],y[3]);
and and1732(ip_27_4,x[27],y[4]);
and and1733(ip_27_5,x[27],y[5]);
and and1734(ip_27_6,x[27],y[6]);
and and1735(ip_27_7,x[27],y[7]);
and and1736(ip_27_8,x[27],y[8]);
and and1737(ip_27_9,x[27],y[9]);
and and1738(ip_27_10,x[27],y[10]);
and and1739(ip_27_11,x[27],y[11]);
and and1740(ip_27_12,x[27],y[12]);
and and1741(ip_27_13,x[27],y[13]);
and and1742(ip_27_14,x[27],y[14]);
and and1743(ip_27_15,x[27],y[15]);
and and1744(ip_27_16,x[27],y[16]);
and and1745(ip_27_17,x[27],y[17]);
and and1746(ip_27_18,x[27],y[18]);
and and1747(ip_27_19,x[27],y[19]);
and and1748(ip_27_20,x[27],y[20]);
and and1749(ip_27_21,x[27],y[21]);
and and1750(ip_27_22,x[27],y[22]);
and and1751(ip_27_23,x[27],y[23]);
and and1752(ip_27_24,x[27],y[24]);
and and1753(ip_27_25,x[27],y[25]);
and and1754(ip_27_26,x[27],y[26]);
and and1755(ip_27_27,x[27],y[27]);
and and1756(ip_27_28,x[27],y[28]);
and and1757(ip_27_29,x[27],y[29]);
and and1758(ip_27_30,x[27],y[30]);
and and1759(ip_27_31,x[27],y[31]);
and and1760(ip_27_32,x[27],y[32]);
and and1761(ip_27_33,x[27],y[33]);
and and1762(ip_27_34,x[27],y[34]);
and and1763(ip_27_35,x[27],y[35]);
and and1764(ip_27_36,x[27],y[36]);
and and1765(ip_27_37,x[27],y[37]);
and and1766(ip_27_38,x[27],y[38]);
and and1767(ip_27_39,x[27],y[39]);
and and1768(ip_27_40,x[27],y[40]);
and and1769(ip_27_41,x[27],y[41]);
and and1770(ip_27_42,x[27],y[42]);
and and1771(ip_27_43,x[27],y[43]);
and and1772(ip_27_44,x[27],y[44]);
and and1773(ip_27_45,x[27],y[45]);
and and1774(ip_27_46,x[27],y[46]);
and and1775(ip_27_47,x[27],y[47]);
and and1776(ip_27_48,x[27],y[48]);
and and1777(ip_27_49,x[27],y[49]);
and and1778(ip_27_50,x[27],y[50]);
and and1779(ip_27_51,x[27],y[51]);
and and1780(ip_27_52,x[27],y[52]);
and and1781(ip_27_53,x[27],y[53]);
and and1782(ip_27_54,x[27],y[54]);
and and1783(ip_27_55,x[27],y[55]);
and and1784(ip_27_56,x[27],y[56]);
and and1785(ip_27_57,x[27],y[57]);
and and1786(ip_27_58,x[27],y[58]);
and and1787(ip_27_59,x[27],y[59]);
and and1788(ip_27_60,x[27],y[60]);
and and1789(ip_27_61,x[27],y[61]);
and and1790(ip_27_62,x[27],y[62]);
and and1791(ip_27_63,x[27],y[63]);
and and1792(ip_28_0,x[28],y[0]);
and and1793(ip_28_1,x[28],y[1]);
and and1794(ip_28_2,x[28],y[2]);
and and1795(ip_28_3,x[28],y[3]);
and and1796(ip_28_4,x[28],y[4]);
and and1797(ip_28_5,x[28],y[5]);
and and1798(ip_28_6,x[28],y[6]);
and and1799(ip_28_7,x[28],y[7]);
and and1800(ip_28_8,x[28],y[8]);
and and1801(ip_28_9,x[28],y[9]);
and and1802(ip_28_10,x[28],y[10]);
and and1803(ip_28_11,x[28],y[11]);
and and1804(ip_28_12,x[28],y[12]);
and and1805(ip_28_13,x[28],y[13]);
and and1806(ip_28_14,x[28],y[14]);
and and1807(ip_28_15,x[28],y[15]);
and and1808(ip_28_16,x[28],y[16]);
and and1809(ip_28_17,x[28],y[17]);
and and1810(ip_28_18,x[28],y[18]);
and and1811(ip_28_19,x[28],y[19]);
and and1812(ip_28_20,x[28],y[20]);
and and1813(ip_28_21,x[28],y[21]);
and and1814(ip_28_22,x[28],y[22]);
and and1815(ip_28_23,x[28],y[23]);
and and1816(ip_28_24,x[28],y[24]);
and and1817(ip_28_25,x[28],y[25]);
and and1818(ip_28_26,x[28],y[26]);
and and1819(ip_28_27,x[28],y[27]);
and and1820(ip_28_28,x[28],y[28]);
and and1821(ip_28_29,x[28],y[29]);
and and1822(ip_28_30,x[28],y[30]);
and and1823(ip_28_31,x[28],y[31]);
and and1824(ip_28_32,x[28],y[32]);
and and1825(ip_28_33,x[28],y[33]);
and and1826(ip_28_34,x[28],y[34]);
and and1827(ip_28_35,x[28],y[35]);
and and1828(ip_28_36,x[28],y[36]);
and and1829(ip_28_37,x[28],y[37]);
and and1830(ip_28_38,x[28],y[38]);
and and1831(ip_28_39,x[28],y[39]);
and and1832(ip_28_40,x[28],y[40]);
and and1833(ip_28_41,x[28],y[41]);
and and1834(ip_28_42,x[28],y[42]);
and and1835(ip_28_43,x[28],y[43]);
and and1836(ip_28_44,x[28],y[44]);
and and1837(ip_28_45,x[28],y[45]);
and and1838(ip_28_46,x[28],y[46]);
and and1839(ip_28_47,x[28],y[47]);
and and1840(ip_28_48,x[28],y[48]);
and and1841(ip_28_49,x[28],y[49]);
and and1842(ip_28_50,x[28],y[50]);
and and1843(ip_28_51,x[28],y[51]);
and and1844(ip_28_52,x[28],y[52]);
and and1845(ip_28_53,x[28],y[53]);
and and1846(ip_28_54,x[28],y[54]);
and and1847(ip_28_55,x[28],y[55]);
and and1848(ip_28_56,x[28],y[56]);
and and1849(ip_28_57,x[28],y[57]);
and and1850(ip_28_58,x[28],y[58]);
and and1851(ip_28_59,x[28],y[59]);
and and1852(ip_28_60,x[28],y[60]);
and and1853(ip_28_61,x[28],y[61]);
and and1854(ip_28_62,x[28],y[62]);
and and1855(ip_28_63,x[28],y[63]);
and and1856(ip_29_0,x[29],y[0]);
and and1857(ip_29_1,x[29],y[1]);
and and1858(ip_29_2,x[29],y[2]);
and and1859(ip_29_3,x[29],y[3]);
and and1860(ip_29_4,x[29],y[4]);
and and1861(ip_29_5,x[29],y[5]);
and and1862(ip_29_6,x[29],y[6]);
and and1863(ip_29_7,x[29],y[7]);
and and1864(ip_29_8,x[29],y[8]);
and and1865(ip_29_9,x[29],y[9]);
and and1866(ip_29_10,x[29],y[10]);
and and1867(ip_29_11,x[29],y[11]);
and and1868(ip_29_12,x[29],y[12]);
and and1869(ip_29_13,x[29],y[13]);
and and1870(ip_29_14,x[29],y[14]);
and and1871(ip_29_15,x[29],y[15]);
and and1872(ip_29_16,x[29],y[16]);
and and1873(ip_29_17,x[29],y[17]);
and and1874(ip_29_18,x[29],y[18]);
and and1875(ip_29_19,x[29],y[19]);
and and1876(ip_29_20,x[29],y[20]);
and and1877(ip_29_21,x[29],y[21]);
and and1878(ip_29_22,x[29],y[22]);
and and1879(ip_29_23,x[29],y[23]);
and and1880(ip_29_24,x[29],y[24]);
and and1881(ip_29_25,x[29],y[25]);
and and1882(ip_29_26,x[29],y[26]);
and and1883(ip_29_27,x[29],y[27]);
and and1884(ip_29_28,x[29],y[28]);
and and1885(ip_29_29,x[29],y[29]);
and and1886(ip_29_30,x[29],y[30]);
and and1887(ip_29_31,x[29],y[31]);
and and1888(ip_29_32,x[29],y[32]);
and and1889(ip_29_33,x[29],y[33]);
and and1890(ip_29_34,x[29],y[34]);
and and1891(ip_29_35,x[29],y[35]);
and and1892(ip_29_36,x[29],y[36]);
and and1893(ip_29_37,x[29],y[37]);
and and1894(ip_29_38,x[29],y[38]);
and and1895(ip_29_39,x[29],y[39]);
and and1896(ip_29_40,x[29],y[40]);
and and1897(ip_29_41,x[29],y[41]);
and and1898(ip_29_42,x[29],y[42]);
and and1899(ip_29_43,x[29],y[43]);
and and1900(ip_29_44,x[29],y[44]);
and and1901(ip_29_45,x[29],y[45]);
and and1902(ip_29_46,x[29],y[46]);
and and1903(ip_29_47,x[29],y[47]);
and and1904(ip_29_48,x[29],y[48]);
and and1905(ip_29_49,x[29],y[49]);
and and1906(ip_29_50,x[29],y[50]);
and and1907(ip_29_51,x[29],y[51]);
and and1908(ip_29_52,x[29],y[52]);
and and1909(ip_29_53,x[29],y[53]);
and and1910(ip_29_54,x[29],y[54]);
and and1911(ip_29_55,x[29],y[55]);
and and1912(ip_29_56,x[29],y[56]);
and and1913(ip_29_57,x[29],y[57]);
and and1914(ip_29_58,x[29],y[58]);
and and1915(ip_29_59,x[29],y[59]);
and and1916(ip_29_60,x[29],y[60]);
and and1917(ip_29_61,x[29],y[61]);
and and1918(ip_29_62,x[29],y[62]);
and and1919(ip_29_63,x[29],y[63]);
and and1920(ip_30_0,x[30],y[0]);
and and1921(ip_30_1,x[30],y[1]);
and and1922(ip_30_2,x[30],y[2]);
and and1923(ip_30_3,x[30],y[3]);
and and1924(ip_30_4,x[30],y[4]);
and and1925(ip_30_5,x[30],y[5]);
and and1926(ip_30_6,x[30],y[6]);
and and1927(ip_30_7,x[30],y[7]);
and and1928(ip_30_8,x[30],y[8]);
and and1929(ip_30_9,x[30],y[9]);
and and1930(ip_30_10,x[30],y[10]);
and and1931(ip_30_11,x[30],y[11]);
and and1932(ip_30_12,x[30],y[12]);
and and1933(ip_30_13,x[30],y[13]);
and and1934(ip_30_14,x[30],y[14]);
and and1935(ip_30_15,x[30],y[15]);
and and1936(ip_30_16,x[30],y[16]);
and and1937(ip_30_17,x[30],y[17]);
and and1938(ip_30_18,x[30],y[18]);
and and1939(ip_30_19,x[30],y[19]);
and and1940(ip_30_20,x[30],y[20]);
and and1941(ip_30_21,x[30],y[21]);
and and1942(ip_30_22,x[30],y[22]);
and and1943(ip_30_23,x[30],y[23]);
and and1944(ip_30_24,x[30],y[24]);
and and1945(ip_30_25,x[30],y[25]);
and and1946(ip_30_26,x[30],y[26]);
and and1947(ip_30_27,x[30],y[27]);
and and1948(ip_30_28,x[30],y[28]);
and and1949(ip_30_29,x[30],y[29]);
and and1950(ip_30_30,x[30],y[30]);
and and1951(ip_30_31,x[30],y[31]);
and and1952(ip_30_32,x[30],y[32]);
and and1953(ip_30_33,x[30],y[33]);
and and1954(ip_30_34,x[30],y[34]);
and and1955(ip_30_35,x[30],y[35]);
and and1956(ip_30_36,x[30],y[36]);
and and1957(ip_30_37,x[30],y[37]);
and and1958(ip_30_38,x[30],y[38]);
and and1959(ip_30_39,x[30],y[39]);
and and1960(ip_30_40,x[30],y[40]);
and and1961(ip_30_41,x[30],y[41]);
and and1962(ip_30_42,x[30],y[42]);
and and1963(ip_30_43,x[30],y[43]);
and and1964(ip_30_44,x[30],y[44]);
and and1965(ip_30_45,x[30],y[45]);
and and1966(ip_30_46,x[30],y[46]);
and and1967(ip_30_47,x[30],y[47]);
and and1968(ip_30_48,x[30],y[48]);
and and1969(ip_30_49,x[30],y[49]);
and and1970(ip_30_50,x[30],y[50]);
and and1971(ip_30_51,x[30],y[51]);
and and1972(ip_30_52,x[30],y[52]);
and and1973(ip_30_53,x[30],y[53]);
and and1974(ip_30_54,x[30],y[54]);
and and1975(ip_30_55,x[30],y[55]);
and and1976(ip_30_56,x[30],y[56]);
and and1977(ip_30_57,x[30],y[57]);
and and1978(ip_30_58,x[30],y[58]);
and and1979(ip_30_59,x[30],y[59]);
and and1980(ip_30_60,x[30],y[60]);
and and1981(ip_30_61,x[30],y[61]);
and and1982(ip_30_62,x[30],y[62]);
and and1983(ip_30_63,x[30],y[63]);
and and1984(ip_31_0,x[31],y[0]);
and and1985(ip_31_1,x[31],y[1]);
and and1986(ip_31_2,x[31],y[2]);
and and1987(ip_31_3,x[31],y[3]);
and and1988(ip_31_4,x[31],y[4]);
and and1989(ip_31_5,x[31],y[5]);
and and1990(ip_31_6,x[31],y[6]);
and and1991(ip_31_7,x[31],y[7]);
and and1992(ip_31_8,x[31],y[8]);
and and1993(ip_31_9,x[31],y[9]);
and and1994(ip_31_10,x[31],y[10]);
and and1995(ip_31_11,x[31],y[11]);
and and1996(ip_31_12,x[31],y[12]);
and and1997(ip_31_13,x[31],y[13]);
and and1998(ip_31_14,x[31],y[14]);
and and1999(ip_31_15,x[31],y[15]);
and and2000(ip_31_16,x[31],y[16]);
and and2001(ip_31_17,x[31],y[17]);
and and2002(ip_31_18,x[31],y[18]);
and and2003(ip_31_19,x[31],y[19]);
and and2004(ip_31_20,x[31],y[20]);
and and2005(ip_31_21,x[31],y[21]);
and and2006(ip_31_22,x[31],y[22]);
and and2007(ip_31_23,x[31],y[23]);
and and2008(ip_31_24,x[31],y[24]);
and and2009(ip_31_25,x[31],y[25]);
and and2010(ip_31_26,x[31],y[26]);
and and2011(ip_31_27,x[31],y[27]);
and and2012(ip_31_28,x[31],y[28]);
and and2013(ip_31_29,x[31],y[29]);
and and2014(ip_31_30,x[31],y[30]);
and and2015(ip_31_31,x[31],y[31]);
and and2016(ip_31_32,x[31],y[32]);
and and2017(ip_31_33,x[31],y[33]);
and and2018(ip_31_34,x[31],y[34]);
and and2019(ip_31_35,x[31],y[35]);
and and2020(ip_31_36,x[31],y[36]);
and and2021(ip_31_37,x[31],y[37]);
and and2022(ip_31_38,x[31],y[38]);
and and2023(ip_31_39,x[31],y[39]);
and and2024(ip_31_40,x[31],y[40]);
and and2025(ip_31_41,x[31],y[41]);
and and2026(ip_31_42,x[31],y[42]);
and and2027(ip_31_43,x[31],y[43]);
and and2028(ip_31_44,x[31],y[44]);
and and2029(ip_31_45,x[31],y[45]);
and and2030(ip_31_46,x[31],y[46]);
and and2031(ip_31_47,x[31],y[47]);
and and2032(ip_31_48,x[31],y[48]);
and and2033(ip_31_49,x[31],y[49]);
and and2034(ip_31_50,x[31],y[50]);
and and2035(ip_31_51,x[31],y[51]);
and and2036(ip_31_52,x[31],y[52]);
and and2037(ip_31_53,x[31],y[53]);
and and2038(ip_31_54,x[31],y[54]);
and and2039(ip_31_55,x[31],y[55]);
and and2040(ip_31_56,x[31],y[56]);
and and2041(ip_31_57,x[31],y[57]);
and and2042(ip_31_58,x[31],y[58]);
and and2043(ip_31_59,x[31],y[59]);
and and2044(ip_31_60,x[31],y[60]);
and and2045(ip_31_61,x[31],y[61]);
and and2046(ip_31_62,x[31],y[62]);
and and2047(ip_31_63,x[31],y[63]);
and and2048(ip_32_0,x[32],y[0]);
and and2049(ip_32_1,x[32],y[1]);
and and2050(ip_32_2,x[32],y[2]);
and and2051(ip_32_3,x[32],y[3]);
and and2052(ip_32_4,x[32],y[4]);
and and2053(ip_32_5,x[32],y[5]);
and and2054(ip_32_6,x[32],y[6]);
and and2055(ip_32_7,x[32],y[7]);
and and2056(ip_32_8,x[32],y[8]);
and and2057(ip_32_9,x[32],y[9]);
and and2058(ip_32_10,x[32],y[10]);
and and2059(ip_32_11,x[32],y[11]);
and and2060(ip_32_12,x[32],y[12]);
and and2061(ip_32_13,x[32],y[13]);
and and2062(ip_32_14,x[32],y[14]);
and and2063(ip_32_15,x[32],y[15]);
and and2064(ip_32_16,x[32],y[16]);
and and2065(ip_32_17,x[32],y[17]);
and and2066(ip_32_18,x[32],y[18]);
and and2067(ip_32_19,x[32],y[19]);
and and2068(ip_32_20,x[32],y[20]);
and and2069(ip_32_21,x[32],y[21]);
and and2070(ip_32_22,x[32],y[22]);
and and2071(ip_32_23,x[32],y[23]);
and and2072(ip_32_24,x[32],y[24]);
and and2073(ip_32_25,x[32],y[25]);
and and2074(ip_32_26,x[32],y[26]);
and and2075(ip_32_27,x[32],y[27]);
and and2076(ip_32_28,x[32],y[28]);
and and2077(ip_32_29,x[32],y[29]);
and and2078(ip_32_30,x[32],y[30]);
and and2079(ip_32_31,x[32],y[31]);
and and2080(ip_32_32,x[32],y[32]);
and and2081(ip_32_33,x[32],y[33]);
and and2082(ip_32_34,x[32],y[34]);
and and2083(ip_32_35,x[32],y[35]);
and and2084(ip_32_36,x[32],y[36]);
and and2085(ip_32_37,x[32],y[37]);
and and2086(ip_32_38,x[32],y[38]);
and and2087(ip_32_39,x[32],y[39]);
and and2088(ip_32_40,x[32],y[40]);
and and2089(ip_32_41,x[32],y[41]);
and and2090(ip_32_42,x[32],y[42]);
and and2091(ip_32_43,x[32],y[43]);
and and2092(ip_32_44,x[32],y[44]);
and and2093(ip_32_45,x[32],y[45]);
and and2094(ip_32_46,x[32],y[46]);
and and2095(ip_32_47,x[32],y[47]);
and and2096(ip_32_48,x[32],y[48]);
and and2097(ip_32_49,x[32],y[49]);
and and2098(ip_32_50,x[32],y[50]);
and and2099(ip_32_51,x[32],y[51]);
and and2100(ip_32_52,x[32],y[52]);
and and2101(ip_32_53,x[32],y[53]);
and and2102(ip_32_54,x[32],y[54]);
and and2103(ip_32_55,x[32],y[55]);
and and2104(ip_32_56,x[32],y[56]);
and and2105(ip_32_57,x[32],y[57]);
and and2106(ip_32_58,x[32],y[58]);
and and2107(ip_32_59,x[32],y[59]);
and and2108(ip_32_60,x[32],y[60]);
and and2109(ip_32_61,x[32],y[61]);
and and2110(ip_32_62,x[32],y[62]);
and and2111(ip_32_63,x[32],y[63]);
and and2112(ip_33_0,x[33],y[0]);
and and2113(ip_33_1,x[33],y[1]);
and and2114(ip_33_2,x[33],y[2]);
and and2115(ip_33_3,x[33],y[3]);
and and2116(ip_33_4,x[33],y[4]);
and and2117(ip_33_5,x[33],y[5]);
and and2118(ip_33_6,x[33],y[6]);
and and2119(ip_33_7,x[33],y[7]);
and and2120(ip_33_8,x[33],y[8]);
and and2121(ip_33_9,x[33],y[9]);
and and2122(ip_33_10,x[33],y[10]);
and and2123(ip_33_11,x[33],y[11]);
and and2124(ip_33_12,x[33],y[12]);
and and2125(ip_33_13,x[33],y[13]);
and and2126(ip_33_14,x[33],y[14]);
and and2127(ip_33_15,x[33],y[15]);
and and2128(ip_33_16,x[33],y[16]);
and and2129(ip_33_17,x[33],y[17]);
and and2130(ip_33_18,x[33],y[18]);
and and2131(ip_33_19,x[33],y[19]);
and and2132(ip_33_20,x[33],y[20]);
and and2133(ip_33_21,x[33],y[21]);
and and2134(ip_33_22,x[33],y[22]);
and and2135(ip_33_23,x[33],y[23]);
and and2136(ip_33_24,x[33],y[24]);
and and2137(ip_33_25,x[33],y[25]);
and and2138(ip_33_26,x[33],y[26]);
and and2139(ip_33_27,x[33],y[27]);
and and2140(ip_33_28,x[33],y[28]);
and and2141(ip_33_29,x[33],y[29]);
and and2142(ip_33_30,x[33],y[30]);
and and2143(ip_33_31,x[33],y[31]);
and and2144(ip_33_32,x[33],y[32]);
and and2145(ip_33_33,x[33],y[33]);
and and2146(ip_33_34,x[33],y[34]);
and and2147(ip_33_35,x[33],y[35]);
and and2148(ip_33_36,x[33],y[36]);
and and2149(ip_33_37,x[33],y[37]);
and and2150(ip_33_38,x[33],y[38]);
and and2151(ip_33_39,x[33],y[39]);
and and2152(ip_33_40,x[33],y[40]);
and and2153(ip_33_41,x[33],y[41]);
and and2154(ip_33_42,x[33],y[42]);
and and2155(ip_33_43,x[33],y[43]);
and and2156(ip_33_44,x[33],y[44]);
and and2157(ip_33_45,x[33],y[45]);
and and2158(ip_33_46,x[33],y[46]);
and and2159(ip_33_47,x[33],y[47]);
and and2160(ip_33_48,x[33],y[48]);
and and2161(ip_33_49,x[33],y[49]);
and and2162(ip_33_50,x[33],y[50]);
and and2163(ip_33_51,x[33],y[51]);
and and2164(ip_33_52,x[33],y[52]);
and and2165(ip_33_53,x[33],y[53]);
and and2166(ip_33_54,x[33],y[54]);
and and2167(ip_33_55,x[33],y[55]);
and and2168(ip_33_56,x[33],y[56]);
and and2169(ip_33_57,x[33],y[57]);
and and2170(ip_33_58,x[33],y[58]);
and and2171(ip_33_59,x[33],y[59]);
and and2172(ip_33_60,x[33],y[60]);
and and2173(ip_33_61,x[33],y[61]);
and and2174(ip_33_62,x[33],y[62]);
and and2175(ip_33_63,x[33],y[63]);
and and2176(ip_34_0,x[34],y[0]);
and and2177(ip_34_1,x[34],y[1]);
and and2178(ip_34_2,x[34],y[2]);
and and2179(ip_34_3,x[34],y[3]);
and and2180(ip_34_4,x[34],y[4]);
and and2181(ip_34_5,x[34],y[5]);
and and2182(ip_34_6,x[34],y[6]);
and and2183(ip_34_7,x[34],y[7]);
and and2184(ip_34_8,x[34],y[8]);
and and2185(ip_34_9,x[34],y[9]);
and and2186(ip_34_10,x[34],y[10]);
and and2187(ip_34_11,x[34],y[11]);
and and2188(ip_34_12,x[34],y[12]);
and and2189(ip_34_13,x[34],y[13]);
and and2190(ip_34_14,x[34],y[14]);
and and2191(ip_34_15,x[34],y[15]);
and and2192(ip_34_16,x[34],y[16]);
and and2193(ip_34_17,x[34],y[17]);
and and2194(ip_34_18,x[34],y[18]);
and and2195(ip_34_19,x[34],y[19]);
and and2196(ip_34_20,x[34],y[20]);
and and2197(ip_34_21,x[34],y[21]);
and and2198(ip_34_22,x[34],y[22]);
and and2199(ip_34_23,x[34],y[23]);
and and2200(ip_34_24,x[34],y[24]);
and and2201(ip_34_25,x[34],y[25]);
and and2202(ip_34_26,x[34],y[26]);
and and2203(ip_34_27,x[34],y[27]);
and and2204(ip_34_28,x[34],y[28]);
and and2205(ip_34_29,x[34],y[29]);
and and2206(ip_34_30,x[34],y[30]);
and and2207(ip_34_31,x[34],y[31]);
and and2208(ip_34_32,x[34],y[32]);
and and2209(ip_34_33,x[34],y[33]);
and and2210(ip_34_34,x[34],y[34]);
and and2211(ip_34_35,x[34],y[35]);
and and2212(ip_34_36,x[34],y[36]);
and and2213(ip_34_37,x[34],y[37]);
and and2214(ip_34_38,x[34],y[38]);
and and2215(ip_34_39,x[34],y[39]);
and and2216(ip_34_40,x[34],y[40]);
and and2217(ip_34_41,x[34],y[41]);
and and2218(ip_34_42,x[34],y[42]);
and and2219(ip_34_43,x[34],y[43]);
and and2220(ip_34_44,x[34],y[44]);
and and2221(ip_34_45,x[34],y[45]);
and and2222(ip_34_46,x[34],y[46]);
and and2223(ip_34_47,x[34],y[47]);
and and2224(ip_34_48,x[34],y[48]);
and and2225(ip_34_49,x[34],y[49]);
and and2226(ip_34_50,x[34],y[50]);
and and2227(ip_34_51,x[34],y[51]);
and and2228(ip_34_52,x[34],y[52]);
and and2229(ip_34_53,x[34],y[53]);
and and2230(ip_34_54,x[34],y[54]);
and and2231(ip_34_55,x[34],y[55]);
and and2232(ip_34_56,x[34],y[56]);
and and2233(ip_34_57,x[34],y[57]);
and and2234(ip_34_58,x[34],y[58]);
and and2235(ip_34_59,x[34],y[59]);
and and2236(ip_34_60,x[34],y[60]);
and and2237(ip_34_61,x[34],y[61]);
and and2238(ip_34_62,x[34],y[62]);
and and2239(ip_34_63,x[34],y[63]);
and and2240(ip_35_0,x[35],y[0]);
and and2241(ip_35_1,x[35],y[1]);
and and2242(ip_35_2,x[35],y[2]);
and and2243(ip_35_3,x[35],y[3]);
and and2244(ip_35_4,x[35],y[4]);
and and2245(ip_35_5,x[35],y[5]);
and and2246(ip_35_6,x[35],y[6]);
and and2247(ip_35_7,x[35],y[7]);
and and2248(ip_35_8,x[35],y[8]);
and and2249(ip_35_9,x[35],y[9]);
and and2250(ip_35_10,x[35],y[10]);
and and2251(ip_35_11,x[35],y[11]);
and and2252(ip_35_12,x[35],y[12]);
and and2253(ip_35_13,x[35],y[13]);
and and2254(ip_35_14,x[35],y[14]);
and and2255(ip_35_15,x[35],y[15]);
and and2256(ip_35_16,x[35],y[16]);
and and2257(ip_35_17,x[35],y[17]);
and and2258(ip_35_18,x[35],y[18]);
and and2259(ip_35_19,x[35],y[19]);
and and2260(ip_35_20,x[35],y[20]);
and and2261(ip_35_21,x[35],y[21]);
and and2262(ip_35_22,x[35],y[22]);
and and2263(ip_35_23,x[35],y[23]);
and and2264(ip_35_24,x[35],y[24]);
and and2265(ip_35_25,x[35],y[25]);
and and2266(ip_35_26,x[35],y[26]);
and and2267(ip_35_27,x[35],y[27]);
and and2268(ip_35_28,x[35],y[28]);
and and2269(ip_35_29,x[35],y[29]);
and and2270(ip_35_30,x[35],y[30]);
and and2271(ip_35_31,x[35],y[31]);
and and2272(ip_35_32,x[35],y[32]);
and and2273(ip_35_33,x[35],y[33]);
and and2274(ip_35_34,x[35],y[34]);
and and2275(ip_35_35,x[35],y[35]);
and and2276(ip_35_36,x[35],y[36]);
and and2277(ip_35_37,x[35],y[37]);
and and2278(ip_35_38,x[35],y[38]);
and and2279(ip_35_39,x[35],y[39]);
and and2280(ip_35_40,x[35],y[40]);
and and2281(ip_35_41,x[35],y[41]);
and and2282(ip_35_42,x[35],y[42]);
and and2283(ip_35_43,x[35],y[43]);
and and2284(ip_35_44,x[35],y[44]);
and and2285(ip_35_45,x[35],y[45]);
and and2286(ip_35_46,x[35],y[46]);
and and2287(ip_35_47,x[35],y[47]);
and and2288(ip_35_48,x[35],y[48]);
and and2289(ip_35_49,x[35],y[49]);
and and2290(ip_35_50,x[35],y[50]);
and and2291(ip_35_51,x[35],y[51]);
and and2292(ip_35_52,x[35],y[52]);
and and2293(ip_35_53,x[35],y[53]);
and and2294(ip_35_54,x[35],y[54]);
and and2295(ip_35_55,x[35],y[55]);
and and2296(ip_35_56,x[35],y[56]);
and and2297(ip_35_57,x[35],y[57]);
and and2298(ip_35_58,x[35],y[58]);
and and2299(ip_35_59,x[35],y[59]);
and and2300(ip_35_60,x[35],y[60]);
and and2301(ip_35_61,x[35],y[61]);
and and2302(ip_35_62,x[35],y[62]);
and and2303(ip_35_63,x[35],y[63]);
and and2304(ip_36_0,x[36],y[0]);
and and2305(ip_36_1,x[36],y[1]);
and and2306(ip_36_2,x[36],y[2]);
and and2307(ip_36_3,x[36],y[3]);
and and2308(ip_36_4,x[36],y[4]);
and and2309(ip_36_5,x[36],y[5]);
and and2310(ip_36_6,x[36],y[6]);
and and2311(ip_36_7,x[36],y[7]);
and and2312(ip_36_8,x[36],y[8]);
and and2313(ip_36_9,x[36],y[9]);
and and2314(ip_36_10,x[36],y[10]);
and and2315(ip_36_11,x[36],y[11]);
and and2316(ip_36_12,x[36],y[12]);
and and2317(ip_36_13,x[36],y[13]);
and and2318(ip_36_14,x[36],y[14]);
and and2319(ip_36_15,x[36],y[15]);
and and2320(ip_36_16,x[36],y[16]);
and and2321(ip_36_17,x[36],y[17]);
and and2322(ip_36_18,x[36],y[18]);
and and2323(ip_36_19,x[36],y[19]);
and and2324(ip_36_20,x[36],y[20]);
and and2325(ip_36_21,x[36],y[21]);
and and2326(ip_36_22,x[36],y[22]);
and and2327(ip_36_23,x[36],y[23]);
and and2328(ip_36_24,x[36],y[24]);
and and2329(ip_36_25,x[36],y[25]);
and and2330(ip_36_26,x[36],y[26]);
and and2331(ip_36_27,x[36],y[27]);
and and2332(ip_36_28,x[36],y[28]);
and and2333(ip_36_29,x[36],y[29]);
and and2334(ip_36_30,x[36],y[30]);
and and2335(ip_36_31,x[36],y[31]);
and and2336(ip_36_32,x[36],y[32]);
and and2337(ip_36_33,x[36],y[33]);
and and2338(ip_36_34,x[36],y[34]);
and and2339(ip_36_35,x[36],y[35]);
and and2340(ip_36_36,x[36],y[36]);
and and2341(ip_36_37,x[36],y[37]);
and and2342(ip_36_38,x[36],y[38]);
and and2343(ip_36_39,x[36],y[39]);
and and2344(ip_36_40,x[36],y[40]);
and and2345(ip_36_41,x[36],y[41]);
and and2346(ip_36_42,x[36],y[42]);
and and2347(ip_36_43,x[36],y[43]);
and and2348(ip_36_44,x[36],y[44]);
and and2349(ip_36_45,x[36],y[45]);
and and2350(ip_36_46,x[36],y[46]);
and and2351(ip_36_47,x[36],y[47]);
and and2352(ip_36_48,x[36],y[48]);
and and2353(ip_36_49,x[36],y[49]);
and and2354(ip_36_50,x[36],y[50]);
and and2355(ip_36_51,x[36],y[51]);
and and2356(ip_36_52,x[36],y[52]);
and and2357(ip_36_53,x[36],y[53]);
and and2358(ip_36_54,x[36],y[54]);
and and2359(ip_36_55,x[36],y[55]);
and and2360(ip_36_56,x[36],y[56]);
and and2361(ip_36_57,x[36],y[57]);
and and2362(ip_36_58,x[36],y[58]);
and and2363(ip_36_59,x[36],y[59]);
and and2364(ip_36_60,x[36],y[60]);
and and2365(ip_36_61,x[36],y[61]);
and and2366(ip_36_62,x[36],y[62]);
and and2367(ip_36_63,x[36],y[63]);
and and2368(ip_37_0,x[37],y[0]);
and and2369(ip_37_1,x[37],y[1]);
and and2370(ip_37_2,x[37],y[2]);
and and2371(ip_37_3,x[37],y[3]);
and and2372(ip_37_4,x[37],y[4]);
and and2373(ip_37_5,x[37],y[5]);
and and2374(ip_37_6,x[37],y[6]);
and and2375(ip_37_7,x[37],y[7]);
and and2376(ip_37_8,x[37],y[8]);
and and2377(ip_37_9,x[37],y[9]);
and and2378(ip_37_10,x[37],y[10]);
and and2379(ip_37_11,x[37],y[11]);
and and2380(ip_37_12,x[37],y[12]);
and and2381(ip_37_13,x[37],y[13]);
and and2382(ip_37_14,x[37],y[14]);
and and2383(ip_37_15,x[37],y[15]);
and and2384(ip_37_16,x[37],y[16]);
and and2385(ip_37_17,x[37],y[17]);
and and2386(ip_37_18,x[37],y[18]);
and and2387(ip_37_19,x[37],y[19]);
and and2388(ip_37_20,x[37],y[20]);
and and2389(ip_37_21,x[37],y[21]);
and and2390(ip_37_22,x[37],y[22]);
and and2391(ip_37_23,x[37],y[23]);
and and2392(ip_37_24,x[37],y[24]);
and and2393(ip_37_25,x[37],y[25]);
and and2394(ip_37_26,x[37],y[26]);
and and2395(ip_37_27,x[37],y[27]);
and and2396(ip_37_28,x[37],y[28]);
and and2397(ip_37_29,x[37],y[29]);
and and2398(ip_37_30,x[37],y[30]);
and and2399(ip_37_31,x[37],y[31]);
and and2400(ip_37_32,x[37],y[32]);
and and2401(ip_37_33,x[37],y[33]);
and and2402(ip_37_34,x[37],y[34]);
and and2403(ip_37_35,x[37],y[35]);
and and2404(ip_37_36,x[37],y[36]);
and and2405(ip_37_37,x[37],y[37]);
and and2406(ip_37_38,x[37],y[38]);
and and2407(ip_37_39,x[37],y[39]);
and and2408(ip_37_40,x[37],y[40]);
and and2409(ip_37_41,x[37],y[41]);
and and2410(ip_37_42,x[37],y[42]);
and and2411(ip_37_43,x[37],y[43]);
and and2412(ip_37_44,x[37],y[44]);
and and2413(ip_37_45,x[37],y[45]);
and and2414(ip_37_46,x[37],y[46]);
and and2415(ip_37_47,x[37],y[47]);
and and2416(ip_37_48,x[37],y[48]);
and and2417(ip_37_49,x[37],y[49]);
and and2418(ip_37_50,x[37],y[50]);
and and2419(ip_37_51,x[37],y[51]);
and and2420(ip_37_52,x[37],y[52]);
and and2421(ip_37_53,x[37],y[53]);
and and2422(ip_37_54,x[37],y[54]);
and and2423(ip_37_55,x[37],y[55]);
and and2424(ip_37_56,x[37],y[56]);
and and2425(ip_37_57,x[37],y[57]);
and and2426(ip_37_58,x[37],y[58]);
and and2427(ip_37_59,x[37],y[59]);
and and2428(ip_37_60,x[37],y[60]);
and and2429(ip_37_61,x[37],y[61]);
and and2430(ip_37_62,x[37],y[62]);
and and2431(ip_37_63,x[37],y[63]);
and and2432(ip_38_0,x[38],y[0]);
and and2433(ip_38_1,x[38],y[1]);
and and2434(ip_38_2,x[38],y[2]);
and and2435(ip_38_3,x[38],y[3]);
and and2436(ip_38_4,x[38],y[4]);
and and2437(ip_38_5,x[38],y[5]);
and and2438(ip_38_6,x[38],y[6]);
and and2439(ip_38_7,x[38],y[7]);
and and2440(ip_38_8,x[38],y[8]);
and and2441(ip_38_9,x[38],y[9]);
and and2442(ip_38_10,x[38],y[10]);
and and2443(ip_38_11,x[38],y[11]);
and and2444(ip_38_12,x[38],y[12]);
and and2445(ip_38_13,x[38],y[13]);
and and2446(ip_38_14,x[38],y[14]);
and and2447(ip_38_15,x[38],y[15]);
and and2448(ip_38_16,x[38],y[16]);
and and2449(ip_38_17,x[38],y[17]);
and and2450(ip_38_18,x[38],y[18]);
and and2451(ip_38_19,x[38],y[19]);
and and2452(ip_38_20,x[38],y[20]);
and and2453(ip_38_21,x[38],y[21]);
and and2454(ip_38_22,x[38],y[22]);
and and2455(ip_38_23,x[38],y[23]);
and and2456(ip_38_24,x[38],y[24]);
and and2457(ip_38_25,x[38],y[25]);
and and2458(ip_38_26,x[38],y[26]);
and and2459(ip_38_27,x[38],y[27]);
and and2460(ip_38_28,x[38],y[28]);
and and2461(ip_38_29,x[38],y[29]);
and and2462(ip_38_30,x[38],y[30]);
and and2463(ip_38_31,x[38],y[31]);
and and2464(ip_38_32,x[38],y[32]);
and and2465(ip_38_33,x[38],y[33]);
and and2466(ip_38_34,x[38],y[34]);
and and2467(ip_38_35,x[38],y[35]);
and and2468(ip_38_36,x[38],y[36]);
and and2469(ip_38_37,x[38],y[37]);
and and2470(ip_38_38,x[38],y[38]);
and and2471(ip_38_39,x[38],y[39]);
and and2472(ip_38_40,x[38],y[40]);
and and2473(ip_38_41,x[38],y[41]);
and and2474(ip_38_42,x[38],y[42]);
and and2475(ip_38_43,x[38],y[43]);
and and2476(ip_38_44,x[38],y[44]);
and and2477(ip_38_45,x[38],y[45]);
and and2478(ip_38_46,x[38],y[46]);
and and2479(ip_38_47,x[38],y[47]);
and and2480(ip_38_48,x[38],y[48]);
and and2481(ip_38_49,x[38],y[49]);
and and2482(ip_38_50,x[38],y[50]);
and and2483(ip_38_51,x[38],y[51]);
and and2484(ip_38_52,x[38],y[52]);
and and2485(ip_38_53,x[38],y[53]);
and and2486(ip_38_54,x[38],y[54]);
and and2487(ip_38_55,x[38],y[55]);
and and2488(ip_38_56,x[38],y[56]);
and and2489(ip_38_57,x[38],y[57]);
and and2490(ip_38_58,x[38],y[58]);
and and2491(ip_38_59,x[38],y[59]);
and and2492(ip_38_60,x[38],y[60]);
and and2493(ip_38_61,x[38],y[61]);
and and2494(ip_38_62,x[38],y[62]);
and and2495(ip_38_63,x[38],y[63]);
and and2496(ip_39_0,x[39],y[0]);
and and2497(ip_39_1,x[39],y[1]);
and and2498(ip_39_2,x[39],y[2]);
and and2499(ip_39_3,x[39],y[3]);
and and2500(ip_39_4,x[39],y[4]);
and and2501(ip_39_5,x[39],y[5]);
and and2502(ip_39_6,x[39],y[6]);
and and2503(ip_39_7,x[39],y[7]);
and and2504(ip_39_8,x[39],y[8]);
and and2505(ip_39_9,x[39],y[9]);
and and2506(ip_39_10,x[39],y[10]);
and and2507(ip_39_11,x[39],y[11]);
and and2508(ip_39_12,x[39],y[12]);
and and2509(ip_39_13,x[39],y[13]);
and and2510(ip_39_14,x[39],y[14]);
and and2511(ip_39_15,x[39],y[15]);
and and2512(ip_39_16,x[39],y[16]);
and and2513(ip_39_17,x[39],y[17]);
and and2514(ip_39_18,x[39],y[18]);
and and2515(ip_39_19,x[39],y[19]);
and and2516(ip_39_20,x[39],y[20]);
and and2517(ip_39_21,x[39],y[21]);
and and2518(ip_39_22,x[39],y[22]);
and and2519(ip_39_23,x[39],y[23]);
and and2520(ip_39_24,x[39],y[24]);
and and2521(ip_39_25,x[39],y[25]);
and and2522(ip_39_26,x[39],y[26]);
and and2523(ip_39_27,x[39],y[27]);
and and2524(ip_39_28,x[39],y[28]);
and and2525(ip_39_29,x[39],y[29]);
and and2526(ip_39_30,x[39],y[30]);
and and2527(ip_39_31,x[39],y[31]);
and and2528(ip_39_32,x[39],y[32]);
and and2529(ip_39_33,x[39],y[33]);
and and2530(ip_39_34,x[39],y[34]);
and and2531(ip_39_35,x[39],y[35]);
and and2532(ip_39_36,x[39],y[36]);
and and2533(ip_39_37,x[39],y[37]);
and and2534(ip_39_38,x[39],y[38]);
and and2535(ip_39_39,x[39],y[39]);
and and2536(ip_39_40,x[39],y[40]);
and and2537(ip_39_41,x[39],y[41]);
and and2538(ip_39_42,x[39],y[42]);
and and2539(ip_39_43,x[39],y[43]);
and and2540(ip_39_44,x[39],y[44]);
and and2541(ip_39_45,x[39],y[45]);
and and2542(ip_39_46,x[39],y[46]);
and and2543(ip_39_47,x[39],y[47]);
and and2544(ip_39_48,x[39],y[48]);
and and2545(ip_39_49,x[39],y[49]);
and and2546(ip_39_50,x[39],y[50]);
and and2547(ip_39_51,x[39],y[51]);
and and2548(ip_39_52,x[39],y[52]);
and and2549(ip_39_53,x[39],y[53]);
and and2550(ip_39_54,x[39],y[54]);
and and2551(ip_39_55,x[39],y[55]);
and and2552(ip_39_56,x[39],y[56]);
and and2553(ip_39_57,x[39],y[57]);
and and2554(ip_39_58,x[39],y[58]);
and and2555(ip_39_59,x[39],y[59]);
and and2556(ip_39_60,x[39],y[60]);
and and2557(ip_39_61,x[39],y[61]);
and and2558(ip_39_62,x[39],y[62]);
and and2559(ip_39_63,x[39],y[63]);
and and2560(ip_40_0,x[40],y[0]);
and and2561(ip_40_1,x[40],y[1]);
and and2562(ip_40_2,x[40],y[2]);
and and2563(ip_40_3,x[40],y[3]);
and and2564(ip_40_4,x[40],y[4]);
and and2565(ip_40_5,x[40],y[5]);
and and2566(ip_40_6,x[40],y[6]);
and and2567(ip_40_7,x[40],y[7]);
and and2568(ip_40_8,x[40],y[8]);
and and2569(ip_40_9,x[40],y[9]);
and and2570(ip_40_10,x[40],y[10]);
and and2571(ip_40_11,x[40],y[11]);
and and2572(ip_40_12,x[40],y[12]);
and and2573(ip_40_13,x[40],y[13]);
and and2574(ip_40_14,x[40],y[14]);
and and2575(ip_40_15,x[40],y[15]);
and and2576(ip_40_16,x[40],y[16]);
and and2577(ip_40_17,x[40],y[17]);
and and2578(ip_40_18,x[40],y[18]);
and and2579(ip_40_19,x[40],y[19]);
and and2580(ip_40_20,x[40],y[20]);
and and2581(ip_40_21,x[40],y[21]);
and and2582(ip_40_22,x[40],y[22]);
and and2583(ip_40_23,x[40],y[23]);
and and2584(ip_40_24,x[40],y[24]);
and and2585(ip_40_25,x[40],y[25]);
and and2586(ip_40_26,x[40],y[26]);
and and2587(ip_40_27,x[40],y[27]);
and and2588(ip_40_28,x[40],y[28]);
and and2589(ip_40_29,x[40],y[29]);
and and2590(ip_40_30,x[40],y[30]);
and and2591(ip_40_31,x[40],y[31]);
and and2592(ip_40_32,x[40],y[32]);
and and2593(ip_40_33,x[40],y[33]);
and and2594(ip_40_34,x[40],y[34]);
and and2595(ip_40_35,x[40],y[35]);
and and2596(ip_40_36,x[40],y[36]);
and and2597(ip_40_37,x[40],y[37]);
and and2598(ip_40_38,x[40],y[38]);
and and2599(ip_40_39,x[40],y[39]);
and and2600(ip_40_40,x[40],y[40]);
and and2601(ip_40_41,x[40],y[41]);
and and2602(ip_40_42,x[40],y[42]);
and and2603(ip_40_43,x[40],y[43]);
and and2604(ip_40_44,x[40],y[44]);
and and2605(ip_40_45,x[40],y[45]);
and and2606(ip_40_46,x[40],y[46]);
and and2607(ip_40_47,x[40],y[47]);
and and2608(ip_40_48,x[40],y[48]);
and and2609(ip_40_49,x[40],y[49]);
and and2610(ip_40_50,x[40],y[50]);
and and2611(ip_40_51,x[40],y[51]);
and and2612(ip_40_52,x[40],y[52]);
and and2613(ip_40_53,x[40],y[53]);
and and2614(ip_40_54,x[40],y[54]);
and and2615(ip_40_55,x[40],y[55]);
and and2616(ip_40_56,x[40],y[56]);
and and2617(ip_40_57,x[40],y[57]);
and and2618(ip_40_58,x[40],y[58]);
and and2619(ip_40_59,x[40],y[59]);
and and2620(ip_40_60,x[40],y[60]);
and and2621(ip_40_61,x[40],y[61]);
and and2622(ip_40_62,x[40],y[62]);
and and2623(ip_40_63,x[40],y[63]);
and and2624(ip_41_0,x[41],y[0]);
and and2625(ip_41_1,x[41],y[1]);
and and2626(ip_41_2,x[41],y[2]);
and and2627(ip_41_3,x[41],y[3]);
and and2628(ip_41_4,x[41],y[4]);
and and2629(ip_41_5,x[41],y[5]);
and and2630(ip_41_6,x[41],y[6]);
and and2631(ip_41_7,x[41],y[7]);
and and2632(ip_41_8,x[41],y[8]);
and and2633(ip_41_9,x[41],y[9]);
and and2634(ip_41_10,x[41],y[10]);
and and2635(ip_41_11,x[41],y[11]);
and and2636(ip_41_12,x[41],y[12]);
and and2637(ip_41_13,x[41],y[13]);
and and2638(ip_41_14,x[41],y[14]);
and and2639(ip_41_15,x[41],y[15]);
and and2640(ip_41_16,x[41],y[16]);
and and2641(ip_41_17,x[41],y[17]);
and and2642(ip_41_18,x[41],y[18]);
and and2643(ip_41_19,x[41],y[19]);
and and2644(ip_41_20,x[41],y[20]);
and and2645(ip_41_21,x[41],y[21]);
and and2646(ip_41_22,x[41],y[22]);
and and2647(ip_41_23,x[41],y[23]);
and and2648(ip_41_24,x[41],y[24]);
and and2649(ip_41_25,x[41],y[25]);
and and2650(ip_41_26,x[41],y[26]);
and and2651(ip_41_27,x[41],y[27]);
and and2652(ip_41_28,x[41],y[28]);
and and2653(ip_41_29,x[41],y[29]);
and and2654(ip_41_30,x[41],y[30]);
and and2655(ip_41_31,x[41],y[31]);
and and2656(ip_41_32,x[41],y[32]);
and and2657(ip_41_33,x[41],y[33]);
and and2658(ip_41_34,x[41],y[34]);
and and2659(ip_41_35,x[41],y[35]);
and and2660(ip_41_36,x[41],y[36]);
and and2661(ip_41_37,x[41],y[37]);
and and2662(ip_41_38,x[41],y[38]);
and and2663(ip_41_39,x[41],y[39]);
and and2664(ip_41_40,x[41],y[40]);
and and2665(ip_41_41,x[41],y[41]);
and and2666(ip_41_42,x[41],y[42]);
and and2667(ip_41_43,x[41],y[43]);
and and2668(ip_41_44,x[41],y[44]);
and and2669(ip_41_45,x[41],y[45]);
and and2670(ip_41_46,x[41],y[46]);
and and2671(ip_41_47,x[41],y[47]);
and and2672(ip_41_48,x[41],y[48]);
and and2673(ip_41_49,x[41],y[49]);
and and2674(ip_41_50,x[41],y[50]);
and and2675(ip_41_51,x[41],y[51]);
and and2676(ip_41_52,x[41],y[52]);
and and2677(ip_41_53,x[41],y[53]);
and and2678(ip_41_54,x[41],y[54]);
and and2679(ip_41_55,x[41],y[55]);
and and2680(ip_41_56,x[41],y[56]);
and and2681(ip_41_57,x[41],y[57]);
and and2682(ip_41_58,x[41],y[58]);
and and2683(ip_41_59,x[41],y[59]);
and and2684(ip_41_60,x[41],y[60]);
and and2685(ip_41_61,x[41],y[61]);
and and2686(ip_41_62,x[41],y[62]);
and and2687(ip_41_63,x[41],y[63]);
and and2688(ip_42_0,x[42],y[0]);
and and2689(ip_42_1,x[42],y[1]);
and and2690(ip_42_2,x[42],y[2]);
and and2691(ip_42_3,x[42],y[3]);
and and2692(ip_42_4,x[42],y[4]);
and and2693(ip_42_5,x[42],y[5]);
and and2694(ip_42_6,x[42],y[6]);
and and2695(ip_42_7,x[42],y[7]);
and and2696(ip_42_8,x[42],y[8]);
and and2697(ip_42_9,x[42],y[9]);
and and2698(ip_42_10,x[42],y[10]);
and and2699(ip_42_11,x[42],y[11]);
and and2700(ip_42_12,x[42],y[12]);
and and2701(ip_42_13,x[42],y[13]);
and and2702(ip_42_14,x[42],y[14]);
and and2703(ip_42_15,x[42],y[15]);
and and2704(ip_42_16,x[42],y[16]);
and and2705(ip_42_17,x[42],y[17]);
and and2706(ip_42_18,x[42],y[18]);
and and2707(ip_42_19,x[42],y[19]);
and and2708(ip_42_20,x[42],y[20]);
and and2709(ip_42_21,x[42],y[21]);
and and2710(ip_42_22,x[42],y[22]);
and and2711(ip_42_23,x[42],y[23]);
and and2712(ip_42_24,x[42],y[24]);
and and2713(ip_42_25,x[42],y[25]);
and and2714(ip_42_26,x[42],y[26]);
and and2715(ip_42_27,x[42],y[27]);
and and2716(ip_42_28,x[42],y[28]);
and and2717(ip_42_29,x[42],y[29]);
and and2718(ip_42_30,x[42],y[30]);
and and2719(ip_42_31,x[42],y[31]);
and and2720(ip_42_32,x[42],y[32]);
and and2721(ip_42_33,x[42],y[33]);
and and2722(ip_42_34,x[42],y[34]);
and and2723(ip_42_35,x[42],y[35]);
and and2724(ip_42_36,x[42],y[36]);
and and2725(ip_42_37,x[42],y[37]);
and and2726(ip_42_38,x[42],y[38]);
and and2727(ip_42_39,x[42],y[39]);
and and2728(ip_42_40,x[42],y[40]);
and and2729(ip_42_41,x[42],y[41]);
and and2730(ip_42_42,x[42],y[42]);
and and2731(ip_42_43,x[42],y[43]);
and and2732(ip_42_44,x[42],y[44]);
and and2733(ip_42_45,x[42],y[45]);
and and2734(ip_42_46,x[42],y[46]);
and and2735(ip_42_47,x[42],y[47]);
and and2736(ip_42_48,x[42],y[48]);
and and2737(ip_42_49,x[42],y[49]);
and and2738(ip_42_50,x[42],y[50]);
and and2739(ip_42_51,x[42],y[51]);
and and2740(ip_42_52,x[42],y[52]);
and and2741(ip_42_53,x[42],y[53]);
and and2742(ip_42_54,x[42],y[54]);
and and2743(ip_42_55,x[42],y[55]);
and and2744(ip_42_56,x[42],y[56]);
and and2745(ip_42_57,x[42],y[57]);
and and2746(ip_42_58,x[42],y[58]);
and and2747(ip_42_59,x[42],y[59]);
and and2748(ip_42_60,x[42],y[60]);
and and2749(ip_42_61,x[42],y[61]);
and and2750(ip_42_62,x[42],y[62]);
and and2751(ip_42_63,x[42],y[63]);
and and2752(ip_43_0,x[43],y[0]);
and and2753(ip_43_1,x[43],y[1]);
and and2754(ip_43_2,x[43],y[2]);
and and2755(ip_43_3,x[43],y[3]);
and and2756(ip_43_4,x[43],y[4]);
and and2757(ip_43_5,x[43],y[5]);
and and2758(ip_43_6,x[43],y[6]);
and and2759(ip_43_7,x[43],y[7]);
and and2760(ip_43_8,x[43],y[8]);
and and2761(ip_43_9,x[43],y[9]);
and and2762(ip_43_10,x[43],y[10]);
and and2763(ip_43_11,x[43],y[11]);
and and2764(ip_43_12,x[43],y[12]);
and and2765(ip_43_13,x[43],y[13]);
and and2766(ip_43_14,x[43],y[14]);
and and2767(ip_43_15,x[43],y[15]);
and and2768(ip_43_16,x[43],y[16]);
and and2769(ip_43_17,x[43],y[17]);
and and2770(ip_43_18,x[43],y[18]);
and and2771(ip_43_19,x[43],y[19]);
and and2772(ip_43_20,x[43],y[20]);
and and2773(ip_43_21,x[43],y[21]);
and and2774(ip_43_22,x[43],y[22]);
and and2775(ip_43_23,x[43],y[23]);
and and2776(ip_43_24,x[43],y[24]);
and and2777(ip_43_25,x[43],y[25]);
and and2778(ip_43_26,x[43],y[26]);
and and2779(ip_43_27,x[43],y[27]);
and and2780(ip_43_28,x[43],y[28]);
and and2781(ip_43_29,x[43],y[29]);
and and2782(ip_43_30,x[43],y[30]);
and and2783(ip_43_31,x[43],y[31]);
and and2784(ip_43_32,x[43],y[32]);
and and2785(ip_43_33,x[43],y[33]);
and and2786(ip_43_34,x[43],y[34]);
and and2787(ip_43_35,x[43],y[35]);
and and2788(ip_43_36,x[43],y[36]);
and and2789(ip_43_37,x[43],y[37]);
and and2790(ip_43_38,x[43],y[38]);
and and2791(ip_43_39,x[43],y[39]);
and and2792(ip_43_40,x[43],y[40]);
and and2793(ip_43_41,x[43],y[41]);
and and2794(ip_43_42,x[43],y[42]);
and and2795(ip_43_43,x[43],y[43]);
and and2796(ip_43_44,x[43],y[44]);
and and2797(ip_43_45,x[43],y[45]);
and and2798(ip_43_46,x[43],y[46]);
and and2799(ip_43_47,x[43],y[47]);
and and2800(ip_43_48,x[43],y[48]);
and and2801(ip_43_49,x[43],y[49]);
and and2802(ip_43_50,x[43],y[50]);
and and2803(ip_43_51,x[43],y[51]);
and and2804(ip_43_52,x[43],y[52]);
and and2805(ip_43_53,x[43],y[53]);
and and2806(ip_43_54,x[43],y[54]);
and and2807(ip_43_55,x[43],y[55]);
and and2808(ip_43_56,x[43],y[56]);
and and2809(ip_43_57,x[43],y[57]);
and and2810(ip_43_58,x[43],y[58]);
and and2811(ip_43_59,x[43],y[59]);
and and2812(ip_43_60,x[43],y[60]);
and and2813(ip_43_61,x[43],y[61]);
and and2814(ip_43_62,x[43],y[62]);
and and2815(ip_43_63,x[43],y[63]);
and and2816(ip_44_0,x[44],y[0]);
and and2817(ip_44_1,x[44],y[1]);
and and2818(ip_44_2,x[44],y[2]);
and and2819(ip_44_3,x[44],y[3]);
and and2820(ip_44_4,x[44],y[4]);
and and2821(ip_44_5,x[44],y[5]);
and and2822(ip_44_6,x[44],y[6]);
and and2823(ip_44_7,x[44],y[7]);
and and2824(ip_44_8,x[44],y[8]);
and and2825(ip_44_9,x[44],y[9]);
and and2826(ip_44_10,x[44],y[10]);
and and2827(ip_44_11,x[44],y[11]);
and and2828(ip_44_12,x[44],y[12]);
and and2829(ip_44_13,x[44],y[13]);
and and2830(ip_44_14,x[44],y[14]);
and and2831(ip_44_15,x[44],y[15]);
and and2832(ip_44_16,x[44],y[16]);
and and2833(ip_44_17,x[44],y[17]);
and and2834(ip_44_18,x[44],y[18]);
and and2835(ip_44_19,x[44],y[19]);
and and2836(ip_44_20,x[44],y[20]);
and and2837(ip_44_21,x[44],y[21]);
and and2838(ip_44_22,x[44],y[22]);
and and2839(ip_44_23,x[44],y[23]);
and and2840(ip_44_24,x[44],y[24]);
and and2841(ip_44_25,x[44],y[25]);
and and2842(ip_44_26,x[44],y[26]);
and and2843(ip_44_27,x[44],y[27]);
and and2844(ip_44_28,x[44],y[28]);
and and2845(ip_44_29,x[44],y[29]);
and and2846(ip_44_30,x[44],y[30]);
and and2847(ip_44_31,x[44],y[31]);
and and2848(ip_44_32,x[44],y[32]);
and and2849(ip_44_33,x[44],y[33]);
and and2850(ip_44_34,x[44],y[34]);
and and2851(ip_44_35,x[44],y[35]);
and and2852(ip_44_36,x[44],y[36]);
and and2853(ip_44_37,x[44],y[37]);
and and2854(ip_44_38,x[44],y[38]);
and and2855(ip_44_39,x[44],y[39]);
and and2856(ip_44_40,x[44],y[40]);
and and2857(ip_44_41,x[44],y[41]);
and and2858(ip_44_42,x[44],y[42]);
and and2859(ip_44_43,x[44],y[43]);
and and2860(ip_44_44,x[44],y[44]);
and and2861(ip_44_45,x[44],y[45]);
and and2862(ip_44_46,x[44],y[46]);
and and2863(ip_44_47,x[44],y[47]);
and and2864(ip_44_48,x[44],y[48]);
and and2865(ip_44_49,x[44],y[49]);
and and2866(ip_44_50,x[44],y[50]);
and and2867(ip_44_51,x[44],y[51]);
and and2868(ip_44_52,x[44],y[52]);
and and2869(ip_44_53,x[44],y[53]);
and and2870(ip_44_54,x[44],y[54]);
and and2871(ip_44_55,x[44],y[55]);
and and2872(ip_44_56,x[44],y[56]);
and and2873(ip_44_57,x[44],y[57]);
and and2874(ip_44_58,x[44],y[58]);
and and2875(ip_44_59,x[44],y[59]);
and and2876(ip_44_60,x[44],y[60]);
and and2877(ip_44_61,x[44],y[61]);
and and2878(ip_44_62,x[44],y[62]);
and and2879(ip_44_63,x[44],y[63]);
and and2880(ip_45_0,x[45],y[0]);
and and2881(ip_45_1,x[45],y[1]);
and and2882(ip_45_2,x[45],y[2]);
and and2883(ip_45_3,x[45],y[3]);
and and2884(ip_45_4,x[45],y[4]);
and and2885(ip_45_5,x[45],y[5]);
and and2886(ip_45_6,x[45],y[6]);
and and2887(ip_45_7,x[45],y[7]);
and and2888(ip_45_8,x[45],y[8]);
and and2889(ip_45_9,x[45],y[9]);
and and2890(ip_45_10,x[45],y[10]);
and and2891(ip_45_11,x[45],y[11]);
and and2892(ip_45_12,x[45],y[12]);
and and2893(ip_45_13,x[45],y[13]);
and and2894(ip_45_14,x[45],y[14]);
and and2895(ip_45_15,x[45],y[15]);
and and2896(ip_45_16,x[45],y[16]);
and and2897(ip_45_17,x[45],y[17]);
and and2898(ip_45_18,x[45],y[18]);
and and2899(ip_45_19,x[45],y[19]);
and and2900(ip_45_20,x[45],y[20]);
and and2901(ip_45_21,x[45],y[21]);
and and2902(ip_45_22,x[45],y[22]);
and and2903(ip_45_23,x[45],y[23]);
and and2904(ip_45_24,x[45],y[24]);
and and2905(ip_45_25,x[45],y[25]);
and and2906(ip_45_26,x[45],y[26]);
and and2907(ip_45_27,x[45],y[27]);
and and2908(ip_45_28,x[45],y[28]);
and and2909(ip_45_29,x[45],y[29]);
and and2910(ip_45_30,x[45],y[30]);
and and2911(ip_45_31,x[45],y[31]);
and and2912(ip_45_32,x[45],y[32]);
and and2913(ip_45_33,x[45],y[33]);
and and2914(ip_45_34,x[45],y[34]);
and and2915(ip_45_35,x[45],y[35]);
and and2916(ip_45_36,x[45],y[36]);
and and2917(ip_45_37,x[45],y[37]);
and and2918(ip_45_38,x[45],y[38]);
and and2919(ip_45_39,x[45],y[39]);
and and2920(ip_45_40,x[45],y[40]);
and and2921(ip_45_41,x[45],y[41]);
and and2922(ip_45_42,x[45],y[42]);
and and2923(ip_45_43,x[45],y[43]);
and and2924(ip_45_44,x[45],y[44]);
and and2925(ip_45_45,x[45],y[45]);
and and2926(ip_45_46,x[45],y[46]);
and and2927(ip_45_47,x[45],y[47]);
and and2928(ip_45_48,x[45],y[48]);
and and2929(ip_45_49,x[45],y[49]);
and and2930(ip_45_50,x[45],y[50]);
and and2931(ip_45_51,x[45],y[51]);
and and2932(ip_45_52,x[45],y[52]);
and and2933(ip_45_53,x[45],y[53]);
and and2934(ip_45_54,x[45],y[54]);
and and2935(ip_45_55,x[45],y[55]);
and and2936(ip_45_56,x[45],y[56]);
and and2937(ip_45_57,x[45],y[57]);
and and2938(ip_45_58,x[45],y[58]);
and and2939(ip_45_59,x[45],y[59]);
and and2940(ip_45_60,x[45],y[60]);
and and2941(ip_45_61,x[45],y[61]);
and and2942(ip_45_62,x[45],y[62]);
and and2943(ip_45_63,x[45],y[63]);
and and2944(ip_46_0,x[46],y[0]);
and and2945(ip_46_1,x[46],y[1]);
and and2946(ip_46_2,x[46],y[2]);
and and2947(ip_46_3,x[46],y[3]);
and and2948(ip_46_4,x[46],y[4]);
and and2949(ip_46_5,x[46],y[5]);
and and2950(ip_46_6,x[46],y[6]);
and and2951(ip_46_7,x[46],y[7]);
and and2952(ip_46_8,x[46],y[8]);
and and2953(ip_46_9,x[46],y[9]);
and and2954(ip_46_10,x[46],y[10]);
and and2955(ip_46_11,x[46],y[11]);
and and2956(ip_46_12,x[46],y[12]);
and and2957(ip_46_13,x[46],y[13]);
and and2958(ip_46_14,x[46],y[14]);
and and2959(ip_46_15,x[46],y[15]);
and and2960(ip_46_16,x[46],y[16]);
and and2961(ip_46_17,x[46],y[17]);
and and2962(ip_46_18,x[46],y[18]);
and and2963(ip_46_19,x[46],y[19]);
and and2964(ip_46_20,x[46],y[20]);
and and2965(ip_46_21,x[46],y[21]);
and and2966(ip_46_22,x[46],y[22]);
and and2967(ip_46_23,x[46],y[23]);
and and2968(ip_46_24,x[46],y[24]);
and and2969(ip_46_25,x[46],y[25]);
and and2970(ip_46_26,x[46],y[26]);
and and2971(ip_46_27,x[46],y[27]);
and and2972(ip_46_28,x[46],y[28]);
and and2973(ip_46_29,x[46],y[29]);
and and2974(ip_46_30,x[46],y[30]);
and and2975(ip_46_31,x[46],y[31]);
and and2976(ip_46_32,x[46],y[32]);
and and2977(ip_46_33,x[46],y[33]);
and and2978(ip_46_34,x[46],y[34]);
and and2979(ip_46_35,x[46],y[35]);
and and2980(ip_46_36,x[46],y[36]);
and and2981(ip_46_37,x[46],y[37]);
and and2982(ip_46_38,x[46],y[38]);
and and2983(ip_46_39,x[46],y[39]);
and and2984(ip_46_40,x[46],y[40]);
and and2985(ip_46_41,x[46],y[41]);
and and2986(ip_46_42,x[46],y[42]);
and and2987(ip_46_43,x[46],y[43]);
and and2988(ip_46_44,x[46],y[44]);
and and2989(ip_46_45,x[46],y[45]);
and and2990(ip_46_46,x[46],y[46]);
and and2991(ip_46_47,x[46],y[47]);
and and2992(ip_46_48,x[46],y[48]);
and and2993(ip_46_49,x[46],y[49]);
and and2994(ip_46_50,x[46],y[50]);
and and2995(ip_46_51,x[46],y[51]);
and and2996(ip_46_52,x[46],y[52]);
and and2997(ip_46_53,x[46],y[53]);
and and2998(ip_46_54,x[46],y[54]);
and and2999(ip_46_55,x[46],y[55]);
and and3000(ip_46_56,x[46],y[56]);
and and3001(ip_46_57,x[46],y[57]);
and and3002(ip_46_58,x[46],y[58]);
and and3003(ip_46_59,x[46],y[59]);
and and3004(ip_46_60,x[46],y[60]);
and and3005(ip_46_61,x[46],y[61]);
and and3006(ip_46_62,x[46],y[62]);
and and3007(ip_46_63,x[46],y[63]);
and and3008(ip_47_0,x[47],y[0]);
and and3009(ip_47_1,x[47],y[1]);
and and3010(ip_47_2,x[47],y[2]);
and and3011(ip_47_3,x[47],y[3]);
and and3012(ip_47_4,x[47],y[4]);
and and3013(ip_47_5,x[47],y[5]);
and and3014(ip_47_6,x[47],y[6]);
and and3015(ip_47_7,x[47],y[7]);
and and3016(ip_47_8,x[47],y[8]);
and and3017(ip_47_9,x[47],y[9]);
and and3018(ip_47_10,x[47],y[10]);
and and3019(ip_47_11,x[47],y[11]);
and and3020(ip_47_12,x[47],y[12]);
and and3021(ip_47_13,x[47],y[13]);
and and3022(ip_47_14,x[47],y[14]);
and and3023(ip_47_15,x[47],y[15]);
and and3024(ip_47_16,x[47],y[16]);
and and3025(ip_47_17,x[47],y[17]);
and and3026(ip_47_18,x[47],y[18]);
and and3027(ip_47_19,x[47],y[19]);
and and3028(ip_47_20,x[47],y[20]);
and and3029(ip_47_21,x[47],y[21]);
and and3030(ip_47_22,x[47],y[22]);
and and3031(ip_47_23,x[47],y[23]);
and and3032(ip_47_24,x[47],y[24]);
and and3033(ip_47_25,x[47],y[25]);
and and3034(ip_47_26,x[47],y[26]);
and and3035(ip_47_27,x[47],y[27]);
and and3036(ip_47_28,x[47],y[28]);
and and3037(ip_47_29,x[47],y[29]);
and and3038(ip_47_30,x[47],y[30]);
and and3039(ip_47_31,x[47],y[31]);
and and3040(ip_47_32,x[47],y[32]);
and and3041(ip_47_33,x[47],y[33]);
and and3042(ip_47_34,x[47],y[34]);
and and3043(ip_47_35,x[47],y[35]);
and and3044(ip_47_36,x[47],y[36]);
and and3045(ip_47_37,x[47],y[37]);
and and3046(ip_47_38,x[47],y[38]);
and and3047(ip_47_39,x[47],y[39]);
and and3048(ip_47_40,x[47],y[40]);
and and3049(ip_47_41,x[47],y[41]);
and and3050(ip_47_42,x[47],y[42]);
and and3051(ip_47_43,x[47],y[43]);
and and3052(ip_47_44,x[47],y[44]);
and and3053(ip_47_45,x[47],y[45]);
and and3054(ip_47_46,x[47],y[46]);
and and3055(ip_47_47,x[47],y[47]);
and and3056(ip_47_48,x[47],y[48]);
and and3057(ip_47_49,x[47],y[49]);
and and3058(ip_47_50,x[47],y[50]);
and and3059(ip_47_51,x[47],y[51]);
and and3060(ip_47_52,x[47],y[52]);
and and3061(ip_47_53,x[47],y[53]);
and and3062(ip_47_54,x[47],y[54]);
and and3063(ip_47_55,x[47],y[55]);
and and3064(ip_47_56,x[47],y[56]);
and and3065(ip_47_57,x[47],y[57]);
and and3066(ip_47_58,x[47],y[58]);
and and3067(ip_47_59,x[47],y[59]);
and and3068(ip_47_60,x[47],y[60]);
and and3069(ip_47_61,x[47],y[61]);
and and3070(ip_47_62,x[47],y[62]);
and and3071(ip_47_63,x[47],y[63]);
and and3072(ip_48_0,x[48],y[0]);
and and3073(ip_48_1,x[48],y[1]);
and and3074(ip_48_2,x[48],y[2]);
and and3075(ip_48_3,x[48],y[3]);
and and3076(ip_48_4,x[48],y[4]);
and and3077(ip_48_5,x[48],y[5]);
and and3078(ip_48_6,x[48],y[6]);
and and3079(ip_48_7,x[48],y[7]);
and and3080(ip_48_8,x[48],y[8]);
and and3081(ip_48_9,x[48],y[9]);
and and3082(ip_48_10,x[48],y[10]);
and and3083(ip_48_11,x[48],y[11]);
and and3084(ip_48_12,x[48],y[12]);
and and3085(ip_48_13,x[48],y[13]);
and and3086(ip_48_14,x[48],y[14]);
and and3087(ip_48_15,x[48],y[15]);
and and3088(ip_48_16,x[48],y[16]);
and and3089(ip_48_17,x[48],y[17]);
and and3090(ip_48_18,x[48],y[18]);
and and3091(ip_48_19,x[48],y[19]);
and and3092(ip_48_20,x[48],y[20]);
and and3093(ip_48_21,x[48],y[21]);
and and3094(ip_48_22,x[48],y[22]);
and and3095(ip_48_23,x[48],y[23]);
and and3096(ip_48_24,x[48],y[24]);
and and3097(ip_48_25,x[48],y[25]);
and and3098(ip_48_26,x[48],y[26]);
and and3099(ip_48_27,x[48],y[27]);
and and3100(ip_48_28,x[48],y[28]);
and and3101(ip_48_29,x[48],y[29]);
and and3102(ip_48_30,x[48],y[30]);
and and3103(ip_48_31,x[48],y[31]);
and and3104(ip_48_32,x[48],y[32]);
and and3105(ip_48_33,x[48],y[33]);
and and3106(ip_48_34,x[48],y[34]);
and and3107(ip_48_35,x[48],y[35]);
and and3108(ip_48_36,x[48],y[36]);
and and3109(ip_48_37,x[48],y[37]);
and and3110(ip_48_38,x[48],y[38]);
and and3111(ip_48_39,x[48],y[39]);
and and3112(ip_48_40,x[48],y[40]);
and and3113(ip_48_41,x[48],y[41]);
and and3114(ip_48_42,x[48],y[42]);
and and3115(ip_48_43,x[48],y[43]);
and and3116(ip_48_44,x[48],y[44]);
and and3117(ip_48_45,x[48],y[45]);
and and3118(ip_48_46,x[48],y[46]);
and and3119(ip_48_47,x[48],y[47]);
and and3120(ip_48_48,x[48],y[48]);
and and3121(ip_48_49,x[48],y[49]);
and and3122(ip_48_50,x[48],y[50]);
and and3123(ip_48_51,x[48],y[51]);
and and3124(ip_48_52,x[48],y[52]);
and and3125(ip_48_53,x[48],y[53]);
and and3126(ip_48_54,x[48],y[54]);
and and3127(ip_48_55,x[48],y[55]);
and and3128(ip_48_56,x[48],y[56]);
and and3129(ip_48_57,x[48],y[57]);
and and3130(ip_48_58,x[48],y[58]);
and and3131(ip_48_59,x[48],y[59]);
and and3132(ip_48_60,x[48],y[60]);
and and3133(ip_48_61,x[48],y[61]);
and and3134(ip_48_62,x[48],y[62]);
and and3135(ip_48_63,x[48],y[63]);
and and3136(ip_49_0,x[49],y[0]);
and and3137(ip_49_1,x[49],y[1]);
and and3138(ip_49_2,x[49],y[2]);
and and3139(ip_49_3,x[49],y[3]);
and and3140(ip_49_4,x[49],y[4]);
and and3141(ip_49_5,x[49],y[5]);
and and3142(ip_49_6,x[49],y[6]);
and and3143(ip_49_7,x[49],y[7]);
and and3144(ip_49_8,x[49],y[8]);
and and3145(ip_49_9,x[49],y[9]);
and and3146(ip_49_10,x[49],y[10]);
and and3147(ip_49_11,x[49],y[11]);
and and3148(ip_49_12,x[49],y[12]);
and and3149(ip_49_13,x[49],y[13]);
and and3150(ip_49_14,x[49],y[14]);
and and3151(ip_49_15,x[49],y[15]);
and and3152(ip_49_16,x[49],y[16]);
and and3153(ip_49_17,x[49],y[17]);
and and3154(ip_49_18,x[49],y[18]);
and and3155(ip_49_19,x[49],y[19]);
and and3156(ip_49_20,x[49],y[20]);
and and3157(ip_49_21,x[49],y[21]);
and and3158(ip_49_22,x[49],y[22]);
and and3159(ip_49_23,x[49],y[23]);
and and3160(ip_49_24,x[49],y[24]);
and and3161(ip_49_25,x[49],y[25]);
and and3162(ip_49_26,x[49],y[26]);
and and3163(ip_49_27,x[49],y[27]);
and and3164(ip_49_28,x[49],y[28]);
and and3165(ip_49_29,x[49],y[29]);
and and3166(ip_49_30,x[49],y[30]);
and and3167(ip_49_31,x[49],y[31]);
and and3168(ip_49_32,x[49],y[32]);
and and3169(ip_49_33,x[49],y[33]);
and and3170(ip_49_34,x[49],y[34]);
and and3171(ip_49_35,x[49],y[35]);
and and3172(ip_49_36,x[49],y[36]);
and and3173(ip_49_37,x[49],y[37]);
and and3174(ip_49_38,x[49],y[38]);
and and3175(ip_49_39,x[49],y[39]);
and and3176(ip_49_40,x[49],y[40]);
and and3177(ip_49_41,x[49],y[41]);
and and3178(ip_49_42,x[49],y[42]);
and and3179(ip_49_43,x[49],y[43]);
and and3180(ip_49_44,x[49],y[44]);
and and3181(ip_49_45,x[49],y[45]);
and and3182(ip_49_46,x[49],y[46]);
and and3183(ip_49_47,x[49],y[47]);
and and3184(ip_49_48,x[49],y[48]);
and and3185(ip_49_49,x[49],y[49]);
and and3186(ip_49_50,x[49],y[50]);
and and3187(ip_49_51,x[49],y[51]);
and and3188(ip_49_52,x[49],y[52]);
and and3189(ip_49_53,x[49],y[53]);
and and3190(ip_49_54,x[49],y[54]);
and and3191(ip_49_55,x[49],y[55]);
and and3192(ip_49_56,x[49],y[56]);
and and3193(ip_49_57,x[49],y[57]);
and and3194(ip_49_58,x[49],y[58]);
and and3195(ip_49_59,x[49],y[59]);
and and3196(ip_49_60,x[49],y[60]);
and and3197(ip_49_61,x[49],y[61]);
and and3198(ip_49_62,x[49],y[62]);
and and3199(ip_49_63,x[49],y[63]);
and and3200(ip_50_0,x[50],y[0]);
and and3201(ip_50_1,x[50],y[1]);
and and3202(ip_50_2,x[50],y[2]);
and and3203(ip_50_3,x[50],y[3]);
and and3204(ip_50_4,x[50],y[4]);
and and3205(ip_50_5,x[50],y[5]);
and and3206(ip_50_6,x[50],y[6]);
and and3207(ip_50_7,x[50],y[7]);
and and3208(ip_50_8,x[50],y[8]);
and and3209(ip_50_9,x[50],y[9]);
and and3210(ip_50_10,x[50],y[10]);
and and3211(ip_50_11,x[50],y[11]);
and and3212(ip_50_12,x[50],y[12]);
and and3213(ip_50_13,x[50],y[13]);
and and3214(ip_50_14,x[50],y[14]);
and and3215(ip_50_15,x[50],y[15]);
and and3216(ip_50_16,x[50],y[16]);
and and3217(ip_50_17,x[50],y[17]);
and and3218(ip_50_18,x[50],y[18]);
and and3219(ip_50_19,x[50],y[19]);
and and3220(ip_50_20,x[50],y[20]);
and and3221(ip_50_21,x[50],y[21]);
and and3222(ip_50_22,x[50],y[22]);
and and3223(ip_50_23,x[50],y[23]);
and and3224(ip_50_24,x[50],y[24]);
and and3225(ip_50_25,x[50],y[25]);
and and3226(ip_50_26,x[50],y[26]);
and and3227(ip_50_27,x[50],y[27]);
and and3228(ip_50_28,x[50],y[28]);
and and3229(ip_50_29,x[50],y[29]);
and and3230(ip_50_30,x[50],y[30]);
and and3231(ip_50_31,x[50],y[31]);
and and3232(ip_50_32,x[50],y[32]);
and and3233(ip_50_33,x[50],y[33]);
and and3234(ip_50_34,x[50],y[34]);
and and3235(ip_50_35,x[50],y[35]);
and and3236(ip_50_36,x[50],y[36]);
and and3237(ip_50_37,x[50],y[37]);
and and3238(ip_50_38,x[50],y[38]);
and and3239(ip_50_39,x[50],y[39]);
and and3240(ip_50_40,x[50],y[40]);
and and3241(ip_50_41,x[50],y[41]);
and and3242(ip_50_42,x[50],y[42]);
and and3243(ip_50_43,x[50],y[43]);
and and3244(ip_50_44,x[50],y[44]);
and and3245(ip_50_45,x[50],y[45]);
and and3246(ip_50_46,x[50],y[46]);
and and3247(ip_50_47,x[50],y[47]);
and and3248(ip_50_48,x[50],y[48]);
and and3249(ip_50_49,x[50],y[49]);
and and3250(ip_50_50,x[50],y[50]);
and and3251(ip_50_51,x[50],y[51]);
and and3252(ip_50_52,x[50],y[52]);
and and3253(ip_50_53,x[50],y[53]);
and and3254(ip_50_54,x[50],y[54]);
and and3255(ip_50_55,x[50],y[55]);
and and3256(ip_50_56,x[50],y[56]);
and and3257(ip_50_57,x[50],y[57]);
and and3258(ip_50_58,x[50],y[58]);
and and3259(ip_50_59,x[50],y[59]);
and and3260(ip_50_60,x[50],y[60]);
and and3261(ip_50_61,x[50],y[61]);
and and3262(ip_50_62,x[50],y[62]);
and and3263(ip_50_63,x[50],y[63]);
and and3264(ip_51_0,x[51],y[0]);
and and3265(ip_51_1,x[51],y[1]);
and and3266(ip_51_2,x[51],y[2]);
and and3267(ip_51_3,x[51],y[3]);
and and3268(ip_51_4,x[51],y[4]);
and and3269(ip_51_5,x[51],y[5]);
and and3270(ip_51_6,x[51],y[6]);
and and3271(ip_51_7,x[51],y[7]);
and and3272(ip_51_8,x[51],y[8]);
and and3273(ip_51_9,x[51],y[9]);
and and3274(ip_51_10,x[51],y[10]);
and and3275(ip_51_11,x[51],y[11]);
and and3276(ip_51_12,x[51],y[12]);
and and3277(ip_51_13,x[51],y[13]);
and and3278(ip_51_14,x[51],y[14]);
and and3279(ip_51_15,x[51],y[15]);
and and3280(ip_51_16,x[51],y[16]);
and and3281(ip_51_17,x[51],y[17]);
and and3282(ip_51_18,x[51],y[18]);
and and3283(ip_51_19,x[51],y[19]);
and and3284(ip_51_20,x[51],y[20]);
and and3285(ip_51_21,x[51],y[21]);
and and3286(ip_51_22,x[51],y[22]);
and and3287(ip_51_23,x[51],y[23]);
and and3288(ip_51_24,x[51],y[24]);
and and3289(ip_51_25,x[51],y[25]);
and and3290(ip_51_26,x[51],y[26]);
and and3291(ip_51_27,x[51],y[27]);
and and3292(ip_51_28,x[51],y[28]);
and and3293(ip_51_29,x[51],y[29]);
and and3294(ip_51_30,x[51],y[30]);
and and3295(ip_51_31,x[51],y[31]);
and and3296(ip_51_32,x[51],y[32]);
and and3297(ip_51_33,x[51],y[33]);
and and3298(ip_51_34,x[51],y[34]);
and and3299(ip_51_35,x[51],y[35]);
and and3300(ip_51_36,x[51],y[36]);
and and3301(ip_51_37,x[51],y[37]);
and and3302(ip_51_38,x[51],y[38]);
and and3303(ip_51_39,x[51],y[39]);
and and3304(ip_51_40,x[51],y[40]);
and and3305(ip_51_41,x[51],y[41]);
and and3306(ip_51_42,x[51],y[42]);
and and3307(ip_51_43,x[51],y[43]);
and and3308(ip_51_44,x[51],y[44]);
and and3309(ip_51_45,x[51],y[45]);
and and3310(ip_51_46,x[51],y[46]);
and and3311(ip_51_47,x[51],y[47]);
and and3312(ip_51_48,x[51],y[48]);
and and3313(ip_51_49,x[51],y[49]);
and and3314(ip_51_50,x[51],y[50]);
and and3315(ip_51_51,x[51],y[51]);
and and3316(ip_51_52,x[51],y[52]);
and and3317(ip_51_53,x[51],y[53]);
and and3318(ip_51_54,x[51],y[54]);
and and3319(ip_51_55,x[51],y[55]);
and and3320(ip_51_56,x[51],y[56]);
and and3321(ip_51_57,x[51],y[57]);
and and3322(ip_51_58,x[51],y[58]);
and and3323(ip_51_59,x[51],y[59]);
and and3324(ip_51_60,x[51],y[60]);
and and3325(ip_51_61,x[51],y[61]);
and and3326(ip_51_62,x[51],y[62]);
and and3327(ip_51_63,x[51],y[63]);
and and3328(ip_52_0,x[52],y[0]);
and and3329(ip_52_1,x[52],y[1]);
and and3330(ip_52_2,x[52],y[2]);
and and3331(ip_52_3,x[52],y[3]);
and and3332(ip_52_4,x[52],y[4]);
and and3333(ip_52_5,x[52],y[5]);
and and3334(ip_52_6,x[52],y[6]);
and and3335(ip_52_7,x[52],y[7]);
and and3336(ip_52_8,x[52],y[8]);
and and3337(ip_52_9,x[52],y[9]);
and and3338(ip_52_10,x[52],y[10]);
and and3339(ip_52_11,x[52],y[11]);
and and3340(ip_52_12,x[52],y[12]);
and and3341(ip_52_13,x[52],y[13]);
and and3342(ip_52_14,x[52],y[14]);
and and3343(ip_52_15,x[52],y[15]);
and and3344(ip_52_16,x[52],y[16]);
and and3345(ip_52_17,x[52],y[17]);
and and3346(ip_52_18,x[52],y[18]);
and and3347(ip_52_19,x[52],y[19]);
and and3348(ip_52_20,x[52],y[20]);
and and3349(ip_52_21,x[52],y[21]);
and and3350(ip_52_22,x[52],y[22]);
and and3351(ip_52_23,x[52],y[23]);
and and3352(ip_52_24,x[52],y[24]);
and and3353(ip_52_25,x[52],y[25]);
and and3354(ip_52_26,x[52],y[26]);
and and3355(ip_52_27,x[52],y[27]);
and and3356(ip_52_28,x[52],y[28]);
and and3357(ip_52_29,x[52],y[29]);
and and3358(ip_52_30,x[52],y[30]);
and and3359(ip_52_31,x[52],y[31]);
and and3360(ip_52_32,x[52],y[32]);
and and3361(ip_52_33,x[52],y[33]);
and and3362(ip_52_34,x[52],y[34]);
and and3363(ip_52_35,x[52],y[35]);
and and3364(ip_52_36,x[52],y[36]);
and and3365(ip_52_37,x[52],y[37]);
and and3366(ip_52_38,x[52],y[38]);
and and3367(ip_52_39,x[52],y[39]);
and and3368(ip_52_40,x[52],y[40]);
and and3369(ip_52_41,x[52],y[41]);
and and3370(ip_52_42,x[52],y[42]);
and and3371(ip_52_43,x[52],y[43]);
and and3372(ip_52_44,x[52],y[44]);
and and3373(ip_52_45,x[52],y[45]);
and and3374(ip_52_46,x[52],y[46]);
and and3375(ip_52_47,x[52],y[47]);
and and3376(ip_52_48,x[52],y[48]);
and and3377(ip_52_49,x[52],y[49]);
and and3378(ip_52_50,x[52],y[50]);
and and3379(ip_52_51,x[52],y[51]);
and and3380(ip_52_52,x[52],y[52]);
and and3381(ip_52_53,x[52],y[53]);
and and3382(ip_52_54,x[52],y[54]);
and and3383(ip_52_55,x[52],y[55]);
and and3384(ip_52_56,x[52],y[56]);
and and3385(ip_52_57,x[52],y[57]);
and and3386(ip_52_58,x[52],y[58]);
and and3387(ip_52_59,x[52],y[59]);
and and3388(ip_52_60,x[52],y[60]);
and and3389(ip_52_61,x[52],y[61]);
and and3390(ip_52_62,x[52],y[62]);
and and3391(ip_52_63,x[52],y[63]);
and and3392(ip_53_0,x[53],y[0]);
and and3393(ip_53_1,x[53],y[1]);
and and3394(ip_53_2,x[53],y[2]);
and and3395(ip_53_3,x[53],y[3]);
and and3396(ip_53_4,x[53],y[4]);
and and3397(ip_53_5,x[53],y[5]);
and and3398(ip_53_6,x[53],y[6]);
and and3399(ip_53_7,x[53],y[7]);
and and3400(ip_53_8,x[53],y[8]);
and and3401(ip_53_9,x[53],y[9]);
and and3402(ip_53_10,x[53],y[10]);
and and3403(ip_53_11,x[53],y[11]);
and and3404(ip_53_12,x[53],y[12]);
and and3405(ip_53_13,x[53],y[13]);
and and3406(ip_53_14,x[53],y[14]);
and and3407(ip_53_15,x[53],y[15]);
and and3408(ip_53_16,x[53],y[16]);
and and3409(ip_53_17,x[53],y[17]);
and and3410(ip_53_18,x[53],y[18]);
and and3411(ip_53_19,x[53],y[19]);
and and3412(ip_53_20,x[53],y[20]);
and and3413(ip_53_21,x[53],y[21]);
and and3414(ip_53_22,x[53],y[22]);
and and3415(ip_53_23,x[53],y[23]);
and and3416(ip_53_24,x[53],y[24]);
and and3417(ip_53_25,x[53],y[25]);
and and3418(ip_53_26,x[53],y[26]);
and and3419(ip_53_27,x[53],y[27]);
and and3420(ip_53_28,x[53],y[28]);
and and3421(ip_53_29,x[53],y[29]);
and and3422(ip_53_30,x[53],y[30]);
and and3423(ip_53_31,x[53],y[31]);
and and3424(ip_53_32,x[53],y[32]);
and and3425(ip_53_33,x[53],y[33]);
and and3426(ip_53_34,x[53],y[34]);
and and3427(ip_53_35,x[53],y[35]);
and and3428(ip_53_36,x[53],y[36]);
and and3429(ip_53_37,x[53],y[37]);
and and3430(ip_53_38,x[53],y[38]);
and and3431(ip_53_39,x[53],y[39]);
and and3432(ip_53_40,x[53],y[40]);
and and3433(ip_53_41,x[53],y[41]);
and and3434(ip_53_42,x[53],y[42]);
and and3435(ip_53_43,x[53],y[43]);
and and3436(ip_53_44,x[53],y[44]);
and and3437(ip_53_45,x[53],y[45]);
and and3438(ip_53_46,x[53],y[46]);
and and3439(ip_53_47,x[53],y[47]);
and and3440(ip_53_48,x[53],y[48]);
and and3441(ip_53_49,x[53],y[49]);
and and3442(ip_53_50,x[53],y[50]);
and and3443(ip_53_51,x[53],y[51]);
and and3444(ip_53_52,x[53],y[52]);
and and3445(ip_53_53,x[53],y[53]);
and and3446(ip_53_54,x[53],y[54]);
and and3447(ip_53_55,x[53],y[55]);
and and3448(ip_53_56,x[53],y[56]);
and and3449(ip_53_57,x[53],y[57]);
and and3450(ip_53_58,x[53],y[58]);
and and3451(ip_53_59,x[53],y[59]);
and and3452(ip_53_60,x[53],y[60]);
and and3453(ip_53_61,x[53],y[61]);
and and3454(ip_53_62,x[53],y[62]);
and and3455(ip_53_63,x[53],y[63]);
and and3456(ip_54_0,x[54],y[0]);
and and3457(ip_54_1,x[54],y[1]);
and and3458(ip_54_2,x[54],y[2]);
and and3459(ip_54_3,x[54],y[3]);
and and3460(ip_54_4,x[54],y[4]);
and and3461(ip_54_5,x[54],y[5]);
and and3462(ip_54_6,x[54],y[6]);
and and3463(ip_54_7,x[54],y[7]);
and and3464(ip_54_8,x[54],y[8]);
and and3465(ip_54_9,x[54],y[9]);
and and3466(ip_54_10,x[54],y[10]);
and and3467(ip_54_11,x[54],y[11]);
and and3468(ip_54_12,x[54],y[12]);
and and3469(ip_54_13,x[54],y[13]);
and and3470(ip_54_14,x[54],y[14]);
and and3471(ip_54_15,x[54],y[15]);
and and3472(ip_54_16,x[54],y[16]);
and and3473(ip_54_17,x[54],y[17]);
and and3474(ip_54_18,x[54],y[18]);
and and3475(ip_54_19,x[54],y[19]);
and and3476(ip_54_20,x[54],y[20]);
and and3477(ip_54_21,x[54],y[21]);
and and3478(ip_54_22,x[54],y[22]);
and and3479(ip_54_23,x[54],y[23]);
and and3480(ip_54_24,x[54],y[24]);
and and3481(ip_54_25,x[54],y[25]);
and and3482(ip_54_26,x[54],y[26]);
and and3483(ip_54_27,x[54],y[27]);
and and3484(ip_54_28,x[54],y[28]);
and and3485(ip_54_29,x[54],y[29]);
and and3486(ip_54_30,x[54],y[30]);
and and3487(ip_54_31,x[54],y[31]);
and and3488(ip_54_32,x[54],y[32]);
and and3489(ip_54_33,x[54],y[33]);
and and3490(ip_54_34,x[54],y[34]);
and and3491(ip_54_35,x[54],y[35]);
and and3492(ip_54_36,x[54],y[36]);
and and3493(ip_54_37,x[54],y[37]);
and and3494(ip_54_38,x[54],y[38]);
and and3495(ip_54_39,x[54],y[39]);
and and3496(ip_54_40,x[54],y[40]);
and and3497(ip_54_41,x[54],y[41]);
and and3498(ip_54_42,x[54],y[42]);
and and3499(ip_54_43,x[54],y[43]);
and and3500(ip_54_44,x[54],y[44]);
and and3501(ip_54_45,x[54],y[45]);
and and3502(ip_54_46,x[54],y[46]);
and and3503(ip_54_47,x[54],y[47]);
and and3504(ip_54_48,x[54],y[48]);
and and3505(ip_54_49,x[54],y[49]);
and and3506(ip_54_50,x[54],y[50]);
and and3507(ip_54_51,x[54],y[51]);
and and3508(ip_54_52,x[54],y[52]);
and and3509(ip_54_53,x[54],y[53]);
and and3510(ip_54_54,x[54],y[54]);
and and3511(ip_54_55,x[54],y[55]);
and and3512(ip_54_56,x[54],y[56]);
and and3513(ip_54_57,x[54],y[57]);
and and3514(ip_54_58,x[54],y[58]);
and and3515(ip_54_59,x[54],y[59]);
and and3516(ip_54_60,x[54],y[60]);
and and3517(ip_54_61,x[54],y[61]);
and and3518(ip_54_62,x[54],y[62]);
and and3519(ip_54_63,x[54],y[63]);
and and3520(ip_55_0,x[55],y[0]);
and and3521(ip_55_1,x[55],y[1]);
and and3522(ip_55_2,x[55],y[2]);
and and3523(ip_55_3,x[55],y[3]);
and and3524(ip_55_4,x[55],y[4]);
and and3525(ip_55_5,x[55],y[5]);
and and3526(ip_55_6,x[55],y[6]);
and and3527(ip_55_7,x[55],y[7]);
and and3528(ip_55_8,x[55],y[8]);
and and3529(ip_55_9,x[55],y[9]);
and and3530(ip_55_10,x[55],y[10]);
and and3531(ip_55_11,x[55],y[11]);
and and3532(ip_55_12,x[55],y[12]);
and and3533(ip_55_13,x[55],y[13]);
and and3534(ip_55_14,x[55],y[14]);
and and3535(ip_55_15,x[55],y[15]);
and and3536(ip_55_16,x[55],y[16]);
and and3537(ip_55_17,x[55],y[17]);
and and3538(ip_55_18,x[55],y[18]);
and and3539(ip_55_19,x[55],y[19]);
and and3540(ip_55_20,x[55],y[20]);
and and3541(ip_55_21,x[55],y[21]);
and and3542(ip_55_22,x[55],y[22]);
and and3543(ip_55_23,x[55],y[23]);
and and3544(ip_55_24,x[55],y[24]);
and and3545(ip_55_25,x[55],y[25]);
and and3546(ip_55_26,x[55],y[26]);
and and3547(ip_55_27,x[55],y[27]);
and and3548(ip_55_28,x[55],y[28]);
and and3549(ip_55_29,x[55],y[29]);
and and3550(ip_55_30,x[55],y[30]);
and and3551(ip_55_31,x[55],y[31]);
and and3552(ip_55_32,x[55],y[32]);
and and3553(ip_55_33,x[55],y[33]);
and and3554(ip_55_34,x[55],y[34]);
and and3555(ip_55_35,x[55],y[35]);
and and3556(ip_55_36,x[55],y[36]);
and and3557(ip_55_37,x[55],y[37]);
and and3558(ip_55_38,x[55],y[38]);
and and3559(ip_55_39,x[55],y[39]);
and and3560(ip_55_40,x[55],y[40]);
and and3561(ip_55_41,x[55],y[41]);
and and3562(ip_55_42,x[55],y[42]);
and and3563(ip_55_43,x[55],y[43]);
and and3564(ip_55_44,x[55],y[44]);
and and3565(ip_55_45,x[55],y[45]);
and and3566(ip_55_46,x[55],y[46]);
and and3567(ip_55_47,x[55],y[47]);
and and3568(ip_55_48,x[55],y[48]);
and and3569(ip_55_49,x[55],y[49]);
and and3570(ip_55_50,x[55],y[50]);
and and3571(ip_55_51,x[55],y[51]);
and and3572(ip_55_52,x[55],y[52]);
and and3573(ip_55_53,x[55],y[53]);
and and3574(ip_55_54,x[55],y[54]);
and and3575(ip_55_55,x[55],y[55]);
and and3576(ip_55_56,x[55],y[56]);
and and3577(ip_55_57,x[55],y[57]);
and and3578(ip_55_58,x[55],y[58]);
and and3579(ip_55_59,x[55],y[59]);
and and3580(ip_55_60,x[55],y[60]);
and and3581(ip_55_61,x[55],y[61]);
and and3582(ip_55_62,x[55],y[62]);
and and3583(ip_55_63,x[55],y[63]);
and and3584(ip_56_0,x[56],y[0]);
and and3585(ip_56_1,x[56],y[1]);
and and3586(ip_56_2,x[56],y[2]);
and and3587(ip_56_3,x[56],y[3]);
and and3588(ip_56_4,x[56],y[4]);
and and3589(ip_56_5,x[56],y[5]);
and and3590(ip_56_6,x[56],y[6]);
and and3591(ip_56_7,x[56],y[7]);
and and3592(ip_56_8,x[56],y[8]);
and and3593(ip_56_9,x[56],y[9]);
and and3594(ip_56_10,x[56],y[10]);
and and3595(ip_56_11,x[56],y[11]);
and and3596(ip_56_12,x[56],y[12]);
and and3597(ip_56_13,x[56],y[13]);
and and3598(ip_56_14,x[56],y[14]);
and and3599(ip_56_15,x[56],y[15]);
and and3600(ip_56_16,x[56],y[16]);
and and3601(ip_56_17,x[56],y[17]);
and and3602(ip_56_18,x[56],y[18]);
and and3603(ip_56_19,x[56],y[19]);
and and3604(ip_56_20,x[56],y[20]);
and and3605(ip_56_21,x[56],y[21]);
and and3606(ip_56_22,x[56],y[22]);
and and3607(ip_56_23,x[56],y[23]);
and and3608(ip_56_24,x[56],y[24]);
and and3609(ip_56_25,x[56],y[25]);
and and3610(ip_56_26,x[56],y[26]);
and and3611(ip_56_27,x[56],y[27]);
and and3612(ip_56_28,x[56],y[28]);
and and3613(ip_56_29,x[56],y[29]);
and and3614(ip_56_30,x[56],y[30]);
and and3615(ip_56_31,x[56],y[31]);
and and3616(ip_56_32,x[56],y[32]);
and and3617(ip_56_33,x[56],y[33]);
and and3618(ip_56_34,x[56],y[34]);
and and3619(ip_56_35,x[56],y[35]);
and and3620(ip_56_36,x[56],y[36]);
and and3621(ip_56_37,x[56],y[37]);
and and3622(ip_56_38,x[56],y[38]);
and and3623(ip_56_39,x[56],y[39]);
and and3624(ip_56_40,x[56],y[40]);
and and3625(ip_56_41,x[56],y[41]);
and and3626(ip_56_42,x[56],y[42]);
and and3627(ip_56_43,x[56],y[43]);
and and3628(ip_56_44,x[56],y[44]);
and and3629(ip_56_45,x[56],y[45]);
and and3630(ip_56_46,x[56],y[46]);
and and3631(ip_56_47,x[56],y[47]);
and and3632(ip_56_48,x[56],y[48]);
and and3633(ip_56_49,x[56],y[49]);
and and3634(ip_56_50,x[56],y[50]);
and and3635(ip_56_51,x[56],y[51]);
and and3636(ip_56_52,x[56],y[52]);
and and3637(ip_56_53,x[56],y[53]);
and and3638(ip_56_54,x[56],y[54]);
and and3639(ip_56_55,x[56],y[55]);
and and3640(ip_56_56,x[56],y[56]);
and and3641(ip_56_57,x[56],y[57]);
and and3642(ip_56_58,x[56],y[58]);
and and3643(ip_56_59,x[56],y[59]);
and and3644(ip_56_60,x[56],y[60]);
and and3645(ip_56_61,x[56],y[61]);
and and3646(ip_56_62,x[56],y[62]);
and and3647(ip_56_63,x[56],y[63]);
and and3648(ip_57_0,x[57],y[0]);
and and3649(ip_57_1,x[57],y[1]);
and and3650(ip_57_2,x[57],y[2]);
and and3651(ip_57_3,x[57],y[3]);
and and3652(ip_57_4,x[57],y[4]);
and and3653(ip_57_5,x[57],y[5]);
and and3654(ip_57_6,x[57],y[6]);
and and3655(ip_57_7,x[57],y[7]);
and and3656(ip_57_8,x[57],y[8]);
and and3657(ip_57_9,x[57],y[9]);
and and3658(ip_57_10,x[57],y[10]);
and and3659(ip_57_11,x[57],y[11]);
and and3660(ip_57_12,x[57],y[12]);
and and3661(ip_57_13,x[57],y[13]);
and and3662(ip_57_14,x[57],y[14]);
and and3663(ip_57_15,x[57],y[15]);
and and3664(ip_57_16,x[57],y[16]);
and and3665(ip_57_17,x[57],y[17]);
and and3666(ip_57_18,x[57],y[18]);
and and3667(ip_57_19,x[57],y[19]);
and and3668(ip_57_20,x[57],y[20]);
and and3669(ip_57_21,x[57],y[21]);
and and3670(ip_57_22,x[57],y[22]);
and and3671(ip_57_23,x[57],y[23]);
and and3672(ip_57_24,x[57],y[24]);
and and3673(ip_57_25,x[57],y[25]);
and and3674(ip_57_26,x[57],y[26]);
and and3675(ip_57_27,x[57],y[27]);
and and3676(ip_57_28,x[57],y[28]);
and and3677(ip_57_29,x[57],y[29]);
and and3678(ip_57_30,x[57],y[30]);
and and3679(ip_57_31,x[57],y[31]);
and and3680(ip_57_32,x[57],y[32]);
and and3681(ip_57_33,x[57],y[33]);
and and3682(ip_57_34,x[57],y[34]);
and and3683(ip_57_35,x[57],y[35]);
and and3684(ip_57_36,x[57],y[36]);
and and3685(ip_57_37,x[57],y[37]);
and and3686(ip_57_38,x[57],y[38]);
and and3687(ip_57_39,x[57],y[39]);
and and3688(ip_57_40,x[57],y[40]);
and and3689(ip_57_41,x[57],y[41]);
and and3690(ip_57_42,x[57],y[42]);
and and3691(ip_57_43,x[57],y[43]);
and and3692(ip_57_44,x[57],y[44]);
and and3693(ip_57_45,x[57],y[45]);
and and3694(ip_57_46,x[57],y[46]);
and and3695(ip_57_47,x[57],y[47]);
and and3696(ip_57_48,x[57],y[48]);
and and3697(ip_57_49,x[57],y[49]);
and and3698(ip_57_50,x[57],y[50]);
and and3699(ip_57_51,x[57],y[51]);
and and3700(ip_57_52,x[57],y[52]);
and and3701(ip_57_53,x[57],y[53]);
and and3702(ip_57_54,x[57],y[54]);
and and3703(ip_57_55,x[57],y[55]);
and and3704(ip_57_56,x[57],y[56]);
and and3705(ip_57_57,x[57],y[57]);
and and3706(ip_57_58,x[57],y[58]);
and and3707(ip_57_59,x[57],y[59]);
and and3708(ip_57_60,x[57],y[60]);
and and3709(ip_57_61,x[57],y[61]);
and and3710(ip_57_62,x[57],y[62]);
and and3711(ip_57_63,x[57],y[63]);
and and3712(ip_58_0,x[58],y[0]);
and and3713(ip_58_1,x[58],y[1]);
and and3714(ip_58_2,x[58],y[2]);
and and3715(ip_58_3,x[58],y[3]);
and and3716(ip_58_4,x[58],y[4]);
and and3717(ip_58_5,x[58],y[5]);
and and3718(ip_58_6,x[58],y[6]);
and and3719(ip_58_7,x[58],y[7]);
and and3720(ip_58_8,x[58],y[8]);
and and3721(ip_58_9,x[58],y[9]);
and and3722(ip_58_10,x[58],y[10]);
and and3723(ip_58_11,x[58],y[11]);
and and3724(ip_58_12,x[58],y[12]);
and and3725(ip_58_13,x[58],y[13]);
and and3726(ip_58_14,x[58],y[14]);
and and3727(ip_58_15,x[58],y[15]);
and and3728(ip_58_16,x[58],y[16]);
and and3729(ip_58_17,x[58],y[17]);
and and3730(ip_58_18,x[58],y[18]);
and and3731(ip_58_19,x[58],y[19]);
and and3732(ip_58_20,x[58],y[20]);
and and3733(ip_58_21,x[58],y[21]);
and and3734(ip_58_22,x[58],y[22]);
and and3735(ip_58_23,x[58],y[23]);
and and3736(ip_58_24,x[58],y[24]);
and and3737(ip_58_25,x[58],y[25]);
and and3738(ip_58_26,x[58],y[26]);
and and3739(ip_58_27,x[58],y[27]);
and and3740(ip_58_28,x[58],y[28]);
and and3741(ip_58_29,x[58],y[29]);
and and3742(ip_58_30,x[58],y[30]);
and and3743(ip_58_31,x[58],y[31]);
and and3744(ip_58_32,x[58],y[32]);
and and3745(ip_58_33,x[58],y[33]);
and and3746(ip_58_34,x[58],y[34]);
and and3747(ip_58_35,x[58],y[35]);
and and3748(ip_58_36,x[58],y[36]);
and and3749(ip_58_37,x[58],y[37]);
and and3750(ip_58_38,x[58],y[38]);
and and3751(ip_58_39,x[58],y[39]);
and and3752(ip_58_40,x[58],y[40]);
and and3753(ip_58_41,x[58],y[41]);
and and3754(ip_58_42,x[58],y[42]);
and and3755(ip_58_43,x[58],y[43]);
and and3756(ip_58_44,x[58],y[44]);
and and3757(ip_58_45,x[58],y[45]);
and and3758(ip_58_46,x[58],y[46]);
and and3759(ip_58_47,x[58],y[47]);
and and3760(ip_58_48,x[58],y[48]);
and and3761(ip_58_49,x[58],y[49]);
and and3762(ip_58_50,x[58],y[50]);
and and3763(ip_58_51,x[58],y[51]);
and and3764(ip_58_52,x[58],y[52]);
and and3765(ip_58_53,x[58],y[53]);
and and3766(ip_58_54,x[58],y[54]);
and and3767(ip_58_55,x[58],y[55]);
and and3768(ip_58_56,x[58],y[56]);
and and3769(ip_58_57,x[58],y[57]);
and and3770(ip_58_58,x[58],y[58]);
and and3771(ip_58_59,x[58],y[59]);
and and3772(ip_58_60,x[58],y[60]);
and and3773(ip_58_61,x[58],y[61]);
and and3774(ip_58_62,x[58],y[62]);
and and3775(ip_58_63,x[58],y[63]);
and and3776(ip_59_0,x[59],y[0]);
and and3777(ip_59_1,x[59],y[1]);
and and3778(ip_59_2,x[59],y[2]);
and and3779(ip_59_3,x[59],y[3]);
and and3780(ip_59_4,x[59],y[4]);
and and3781(ip_59_5,x[59],y[5]);
and and3782(ip_59_6,x[59],y[6]);
and and3783(ip_59_7,x[59],y[7]);
and and3784(ip_59_8,x[59],y[8]);
and and3785(ip_59_9,x[59],y[9]);
and and3786(ip_59_10,x[59],y[10]);
and and3787(ip_59_11,x[59],y[11]);
and and3788(ip_59_12,x[59],y[12]);
and and3789(ip_59_13,x[59],y[13]);
and and3790(ip_59_14,x[59],y[14]);
and and3791(ip_59_15,x[59],y[15]);
and and3792(ip_59_16,x[59],y[16]);
and and3793(ip_59_17,x[59],y[17]);
and and3794(ip_59_18,x[59],y[18]);
and and3795(ip_59_19,x[59],y[19]);
and and3796(ip_59_20,x[59],y[20]);
and and3797(ip_59_21,x[59],y[21]);
and and3798(ip_59_22,x[59],y[22]);
and and3799(ip_59_23,x[59],y[23]);
and and3800(ip_59_24,x[59],y[24]);
and and3801(ip_59_25,x[59],y[25]);
and and3802(ip_59_26,x[59],y[26]);
and and3803(ip_59_27,x[59],y[27]);
and and3804(ip_59_28,x[59],y[28]);
and and3805(ip_59_29,x[59],y[29]);
and and3806(ip_59_30,x[59],y[30]);
and and3807(ip_59_31,x[59],y[31]);
and and3808(ip_59_32,x[59],y[32]);
and and3809(ip_59_33,x[59],y[33]);
and and3810(ip_59_34,x[59],y[34]);
and and3811(ip_59_35,x[59],y[35]);
and and3812(ip_59_36,x[59],y[36]);
and and3813(ip_59_37,x[59],y[37]);
and and3814(ip_59_38,x[59],y[38]);
and and3815(ip_59_39,x[59],y[39]);
and and3816(ip_59_40,x[59],y[40]);
and and3817(ip_59_41,x[59],y[41]);
and and3818(ip_59_42,x[59],y[42]);
and and3819(ip_59_43,x[59],y[43]);
and and3820(ip_59_44,x[59],y[44]);
and and3821(ip_59_45,x[59],y[45]);
and and3822(ip_59_46,x[59],y[46]);
and and3823(ip_59_47,x[59],y[47]);
and and3824(ip_59_48,x[59],y[48]);
and and3825(ip_59_49,x[59],y[49]);
and and3826(ip_59_50,x[59],y[50]);
and and3827(ip_59_51,x[59],y[51]);
and and3828(ip_59_52,x[59],y[52]);
and and3829(ip_59_53,x[59],y[53]);
and and3830(ip_59_54,x[59],y[54]);
and and3831(ip_59_55,x[59],y[55]);
and and3832(ip_59_56,x[59],y[56]);
and and3833(ip_59_57,x[59],y[57]);
and and3834(ip_59_58,x[59],y[58]);
and and3835(ip_59_59,x[59],y[59]);
and and3836(ip_59_60,x[59],y[60]);
and and3837(ip_59_61,x[59],y[61]);
and and3838(ip_59_62,x[59],y[62]);
and and3839(ip_59_63,x[59],y[63]);
and and3840(ip_60_0,x[60],y[0]);
and and3841(ip_60_1,x[60],y[1]);
and and3842(ip_60_2,x[60],y[2]);
and and3843(ip_60_3,x[60],y[3]);
and and3844(ip_60_4,x[60],y[4]);
and and3845(ip_60_5,x[60],y[5]);
and and3846(ip_60_6,x[60],y[6]);
and and3847(ip_60_7,x[60],y[7]);
and and3848(ip_60_8,x[60],y[8]);
and and3849(ip_60_9,x[60],y[9]);
and and3850(ip_60_10,x[60],y[10]);
and and3851(ip_60_11,x[60],y[11]);
and and3852(ip_60_12,x[60],y[12]);
and and3853(ip_60_13,x[60],y[13]);
and and3854(ip_60_14,x[60],y[14]);
and and3855(ip_60_15,x[60],y[15]);
and and3856(ip_60_16,x[60],y[16]);
and and3857(ip_60_17,x[60],y[17]);
and and3858(ip_60_18,x[60],y[18]);
and and3859(ip_60_19,x[60],y[19]);
and and3860(ip_60_20,x[60],y[20]);
and and3861(ip_60_21,x[60],y[21]);
and and3862(ip_60_22,x[60],y[22]);
and and3863(ip_60_23,x[60],y[23]);
and and3864(ip_60_24,x[60],y[24]);
and and3865(ip_60_25,x[60],y[25]);
and and3866(ip_60_26,x[60],y[26]);
and and3867(ip_60_27,x[60],y[27]);
and and3868(ip_60_28,x[60],y[28]);
and and3869(ip_60_29,x[60],y[29]);
and and3870(ip_60_30,x[60],y[30]);
and and3871(ip_60_31,x[60],y[31]);
and and3872(ip_60_32,x[60],y[32]);
and and3873(ip_60_33,x[60],y[33]);
and and3874(ip_60_34,x[60],y[34]);
and and3875(ip_60_35,x[60],y[35]);
and and3876(ip_60_36,x[60],y[36]);
and and3877(ip_60_37,x[60],y[37]);
and and3878(ip_60_38,x[60],y[38]);
and and3879(ip_60_39,x[60],y[39]);
and and3880(ip_60_40,x[60],y[40]);
and and3881(ip_60_41,x[60],y[41]);
and and3882(ip_60_42,x[60],y[42]);
and and3883(ip_60_43,x[60],y[43]);
and and3884(ip_60_44,x[60],y[44]);
and and3885(ip_60_45,x[60],y[45]);
and and3886(ip_60_46,x[60],y[46]);
and and3887(ip_60_47,x[60],y[47]);
and and3888(ip_60_48,x[60],y[48]);
and and3889(ip_60_49,x[60],y[49]);
and and3890(ip_60_50,x[60],y[50]);
and and3891(ip_60_51,x[60],y[51]);
and and3892(ip_60_52,x[60],y[52]);
and and3893(ip_60_53,x[60],y[53]);
and and3894(ip_60_54,x[60],y[54]);
and and3895(ip_60_55,x[60],y[55]);
and and3896(ip_60_56,x[60],y[56]);
and and3897(ip_60_57,x[60],y[57]);
and and3898(ip_60_58,x[60],y[58]);
and and3899(ip_60_59,x[60],y[59]);
and and3900(ip_60_60,x[60],y[60]);
and and3901(ip_60_61,x[60],y[61]);
and and3902(ip_60_62,x[60],y[62]);
and and3903(ip_60_63,x[60],y[63]);
and and3904(ip_61_0,x[61],y[0]);
and and3905(ip_61_1,x[61],y[1]);
and and3906(ip_61_2,x[61],y[2]);
and and3907(ip_61_3,x[61],y[3]);
and and3908(ip_61_4,x[61],y[4]);
and and3909(ip_61_5,x[61],y[5]);
and and3910(ip_61_6,x[61],y[6]);
and and3911(ip_61_7,x[61],y[7]);
and and3912(ip_61_8,x[61],y[8]);
and and3913(ip_61_9,x[61],y[9]);
and and3914(ip_61_10,x[61],y[10]);
and and3915(ip_61_11,x[61],y[11]);
and and3916(ip_61_12,x[61],y[12]);
and and3917(ip_61_13,x[61],y[13]);
and and3918(ip_61_14,x[61],y[14]);
and and3919(ip_61_15,x[61],y[15]);
and and3920(ip_61_16,x[61],y[16]);
and and3921(ip_61_17,x[61],y[17]);
and and3922(ip_61_18,x[61],y[18]);
and and3923(ip_61_19,x[61],y[19]);
and and3924(ip_61_20,x[61],y[20]);
and and3925(ip_61_21,x[61],y[21]);
and and3926(ip_61_22,x[61],y[22]);
and and3927(ip_61_23,x[61],y[23]);
and and3928(ip_61_24,x[61],y[24]);
and and3929(ip_61_25,x[61],y[25]);
and and3930(ip_61_26,x[61],y[26]);
and and3931(ip_61_27,x[61],y[27]);
and and3932(ip_61_28,x[61],y[28]);
and and3933(ip_61_29,x[61],y[29]);
and and3934(ip_61_30,x[61],y[30]);
and and3935(ip_61_31,x[61],y[31]);
and and3936(ip_61_32,x[61],y[32]);
and and3937(ip_61_33,x[61],y[33]);
and and3938(ip_61_34,x[61],y[34]);
and and3939(ip_61_35,x[61],y[35]);
and and3940(ip_61_36,x[61],y[36]);
and and3941(ip_61_37,x[61],y[37]);
and and3942(ip_61_38,x[61],y[38]);
and and3943(ip_61_39,x[61],y[39]);
and and3944(ip_61_40,x[61],y[40]);
and and3945(ip_61_41,x[61],y[41]);
and and3946(ip_61_42,x[61],y[42]);
and and3947(ip_61_43,x[61],y[43]);
and and3948(ip_61_44,x[61],y[44]);
and and3949(ip_61_45,x[61],y[45]);
and and3950(ip_61_46,x[61],y[46]);
and and3951(ip_61_47,x[61],y[47]);
and and3952(ip_61_48,x[61],y[48]);
and and3953(ip_61_49,x[61],y[49]);
and and3954(ip_61_50,x[61],y[50]);
and and3955(ip_61_51,x[61],y[51]);
and and3956(ip_61_52,x[61],y[52]);
and and3957(ip_61_53,x[61],y[53]);
and and3958(ip_61_54,x[61],y[54]);
and and3959(ip_61_55,x[61],y[55]);
and and3960(ip_61_56,x[61],y[56]);
and and3961(ip_61_57,x[61],y[57]);
and and3962(ip_61_58,x[61],y[58]);
and and3963(ip_61_59,x[61],y[59]);
and and3964(ip_61_60,x[61],y[60]);
and and3965(ip_61_61,x[61],y[61]);
and and3966(ip_61_62,x[61],y[62]);
and and3967(ip_61_63,x[61],y[63]);
and and3968(ip_62_0,x[62],y[0]);
and and3969(ip_62_1,x[62],y[1]);
and and3970(ip_62_2,x[62],y[2]);
and and3971(ip_62_3,x[62],y[3]);
and and3972(ip_62_4,x[62],y[4]);
and and3973(ip_62_5,x[62],y[5]);
and and3974(ip_62_6,x[62],y[6]);
and and3975(ip_62_7,x[62],y[7]);
and and3976(ip_62_8,x[62],y[8]);
and and3977(ip_62_9,x[62],y[9]);
and and3978(ip_62_10,x[62],y[10]);
and and3979(ip_62_11,x[62],y[11]);
and and3980(ip_62_12,x[62],y[12]);
and and3981(ip_62_13,x[62],y[13]);
and and3982(ip_62_14,x[62],y[14]);
and and3983(ip_62_15,x[62],y[15]);
and and3984(ip_62_16,x[62],y[16]);
and and3985(ip_62_17,x[62],y[17]);
and and3986(ip_62_18,x[62],y[18]);
and and3987(ip_62_19,x[62],y[19]);
and and3988(ip_62_20,x[62],y[20]);
and and3989(ip_62_21,x[62],y[21]);
and and3990(ip_62_22,x[62],y[22]);
and and3991(ip_62_23,x[62],y[23]);
and and3992(ip_62_24,x[62],y[24]);
and and3993(ip_62_25,x[62],y[25]);
and and3994(ip_62_26,x[62],y[26]);
and and3995(ip_62_27,x[62],y[27]);
and and3996(ip_62_28,x[62],y[28]);
and and3997(ip_62_29,x[62],y[29]);
and and3998(ip_62_30,x[62],y[30]);
and and3999(ip_62_31,x[62],y[31]);
and and4000(ip_62_32,x[62],y[32]);
and and4001(ip_62_33,x[62],y[33]);
and and4002(ip_62_34,x[62],y[34]);
and and4003(ip_62_35,x[62],y[35]);
and and4004(ip_62_36,x[62],y[36]);
and and4005(ip_62_37,x[62],y[37]);
and and4006(ip_62_38,x[62],y[38]);
and and4007(ip_62_39,x[62],y[39]);
and and4008(ip_62_40,x[62],y[40]);
and and4009(ip_62_41,x[62],y[41]);
and and4010(ip_62_42,x[62],y[42]);
and and4011(ip_62_43,x[62],y[43]);
and and4012(ip_62_44,x[62],y[44]);
and and4013(ip_62_45,x[62],y[45]);
and and4014(ip_62_46,x[62],y[46]);
and and4015(ip_62_47,x[62],y[47]);
and and4016(ip_62_48,x[62],y[48]);
and and4017(ip_62_49,x[62],y[49]);
and and4018(ip_62_50,x[62],y[50]);
and and4019(ip_62_51,x[62],y[51]);
and and4020(ip_62_52,x[62],y[52]);
and and4021(ip_62_53,x[62],y[53]);
and and4022(ip_62_54,x[62],y[54]);
and and4023(ip_62_55,x[62],y[55]);
and and4024(ip_62_56,x[62],y[56]);
and and4025(ip_62_57,x[62],y[57]);
and and4026(ip_62_58,x[62],y[58]);
and and4027(ip_62_59,x[62],y[59]);
and and4028(ip_62_60,x[62],y[60]);
and and4029(ip_62_61,x[62],y[61]);
and and4030(ip_62_62,x[62],y[62]);
and and4031(ip_62_63,x[62],y[63]);
and and4032(ip_63_0,x[63],y[0]);
and and4033(ip_63_1,x[63],y[1]);
and and4034(ip_63_2,x[63],y[2]);
and and4035(ip_63_3,x[63],y[3]);
and and4036(ip_63_4,x[63],y[4]);
and and4037(ip_63_5,x[63],y[5]);
and and4038(ip_63_6,x[63],y[6]);
and and4039(ip_63_7,x[63],y[7]);
and and4040(ip_63_8,x[63],y[8]);
and and4041(ip_63_9,x[63],y[9]);
and and4042(ip_63_10,x[63],y[10]);
and and4043(ip_63_11,x[63],y[11]);
and and4044(ip_63_12,x[63],y[12]);
and and4045(ip_63_13,x[63],y[13]);
and and4046(ip_63_14,x[63],y[14]);
and and4047(ip_63_15,x[63],y[15]);
and and4048(ip_63_16,x[63],y[16]);
and and4049(ip_63_17,x[63],y[17]);
and and4050(ip_63_18,x[63],y[18]);
and and4051(ip_63_19,x[63],y[19]);
and and4052(ip_63_20,x[63],y[20]);
and and4053(ip_63_21,x[63],y[21]);
and and4054(ip_63_22,x[63],y[22]);
and and4055(ip_63_23,x[63],y[23]);
and and4056(ip_63_24,x[63],y[24]);
and and4057(ip_63_25,x[63],y[25]);
and and4058(ip_63_26,x[63],y[26]);
and and4059(ip_63_27,x[63],y[27]);
and and4060(ip_63_28,x[63],y[28]);
and and4061(ip_63_29,x[63],y[29]);
and and4062(ip_63_30,x[63],y[30]);
and and4063(ip_63_31,x[63],y[31]);
and and4064(ip_63_32,x[63],y[32]);
and and4065(ip_63_33,x[63],y[33]);
and and4066(ip_63_34,x[63],y[34]);
and and4067(ip_63_35,x[63],y[35]);
and and4068(ip_63_36,x[63],y[36]);
and and4069(ip_63_37,x[63],y[37]);
and and4070(ip_63_38,x[63],y[38]);
and and4071(ip_63_39,x[63],y[39]);
and and4072(ip_63_40,x[63],y[40]);
and and4073(ip_63_41,x[63],y[41]);
and and4074(ip_63_42,x[63],y[42]);
and and4075(ip_63_43,x[63],y[43]);
and and4076(ip_63_44,x[63],y[44]);
and and4077(ip_63_45,x[63],y[45]);
and and4078(ip_63_46,x[63],y[46]);
and and4079(ip_63_47,x[63],y[47]);
and and4080(ip_63_48,x[63],y[48]);
and and4081(ip_63_49,x[63],y[49]);
and and4082(ip_63_50,x[63],y[50]);
and and4083(ip_63_51,x[63],y[51]);
and and4084(ip_63_52,x[63],y[52]);
and and4085(ip_63_53,x[63],y[53]);
and and4086(ip_63_54,x[63],y[54]);
and and4087(ip_63_55,x[63],y[55]);
and and4088(ip_63_56,x[63],y[56]);
and and4089(ip_63_57,x[63],y[57]);
and and4090(ip_63_58,x[63],y[58]);
and and4091(ip_63_59,x[63],y[59]);
and and4092(ip_63_60,x[63],y[60]);
and and4093(ip_63_61,x[63],y[61]);
and and4094(ip_63_62,x[63],y[62]);
and and4095(ip_63_63,x[63],y[63]);
HA ha0(ip_0_2,ip_1_1,p0,p1);
FA fa0(ip_0_3,ip_1_2,ip_2_1,p2,p3);
HA ha1(ip_3_0,p0,p4,p5);
FA fa1(ip_0_4,ip_1_3,ip_2_2,p6,p7);
HA ha2(ip_3_1,ip_4_0,p8,p9);
FA fa2(p9,p4,p7,p10,p11);
FA fa3(ip_0_5,ip_1_4,ip_2_3,p12,p13);
HA ha3(ip_3_2,ip_4_1,p14,p15);
FA fa4(ip_5_0,p15,p8,p16,p17);
FA fa5(p13,p17,p6,p18,p19);
HA ha4(ip_0_6,ip_1_5,p20,p21);
FA fa6(ip_2_4,ip_3_3,ip_4_2,p22,p23);
FA fa7(ip_5_1,ip_6_0,p14,p24,p25);
FA fa8(p21,p23,p25,p26,p27);
FA fa9(p12,p16,p27,p28,p29);
HA ha5(ip_0_7,ip_1_6,p30,p31);
HA ha6(ip_2_5,ip_3_4,p32,p33);
FA fa10(ip_4_3,ip_5_2,ip_6_1,p34,p35);
FA fa11(ip_7_0,p20,p31,p36,p37);
HA ha7(p33,p35,p38,p39);
FA fa12(p22,p24,p37,p40,p41);
FA fa13(p39,p26,p41,p42,p43);
FA fa14(ip_0_8,ip_1_7,ip_2_6,p44,p45);
FA fa15(ip_3_5,ip_4_4,ip_5_3,p46,p47);
FA fa16(ip_6_2,ip_7_1,ip_8_0,p48,p49);
FA fa17(p30,p32,p45,p50,p51);
FA fa18(p47,p49,p34,p52,p53);
FA fa19(p38,p51,p36,p54,p55);
HA ha8(p53,p55,p56,p57);
FA fa20(p40,p57,p42,p58,p59);
FA fa21(ip_0_9,ip_1_8,ip_2_7,p60,p61);
HA ha9(ip_3_6,ip_4_5,p62,p63);
FA fa22(ip_5_4,ip_6_3,ip_7_2,p64,p65);
FA fa23(ip_8_1,ip_9_0,p63,p66,p67);
HA ha10(p61,p65,p68,p69);
FA fa24(p67,p44,p46,p70,p71);
FA fa25(p48,p69,p50,p72,p73);
FA fa26(p52,p71,p73,p74,p75);
FA fa27(p54,p56,p75,p76,p77);
FA fa28(ip_0_10,ip_1_9,ip_2_8,p78,p79);
HA ha11(ip_3_7,ip_4_6,p80,p81);
FA fa29(ip_5_5,ip_6_4,ip_7_3,p82,p83);
HA ha12(ip_8_2,ip_9_1,p84,p85);
FA fa30(ip_10_0,p62,p81,p86,p87);
FA fa31(p85,p79,p83,p88,p89);
FA fa32(p60,p64,p66,p90,p91);
FA fa33(p68,p87,p89,p92,p93);
FA fa34(p91,p93,p70,p94,p95);
HA ha13(p72,p95,p96,p97);
FA fa35(p74,p97,p76,p98,p99);
FA fa36(ip_0_11,ip_1_10,ip_2_9,p100,p101);
FA fa37(ip_3_8,ip_4_7,ip_5_6,p102,p103);
FA fa38(ip_6_5,ip_7_4,ip_8_3,p104,p105);
FA fa39(ip_9_2,ip_10_1,ip_11_0,p106,p107);
HA ha14(p80,p84,p108,p109);
FA fa40(p101,p103,p105,p110,p111);
HA ha15(p107,p109,p112,p113);
FA fa41(p113,p78,p82,p114,p115);
HA ha16(p111,p86,p116,p117);
HA ha17(p115,p117,p118,p119);
FA fa42(p88,p119,p90,p120,p121);
FA fa43(p92,p121,p94,p122,p123);
FA fa44(p96,p123,p98,p124,p125);
HA ha18(ip_0_12,ip_1_11,p126,p127);
FA fa45(ip_2_10,ip_3_9,ip_4_8,p128,p129);
FA fa46(ip_5_7,ip_6_6,ip_7_5,p130,p131);
HA ha19(ip_8_4,ip_9_3,p132,p133);
FA fa47(ip_10_2,ip_11_1,ip_12_0,p134,p135);
FA fa48(p127,p133,p108,p136,p137);
FA fa49(p129,p131,p135,p138,p139);
HA ha20(p100,p102,p140,p141);
FA fa50(p104,p106,p112,p142,p143);
FA fa51(p137,p139,p141,p144,p145);
HA ha21(p110,p116,p146,p147);
FA fa52(p143,p114,p118,p148,p149);
FA fa53(p145,p147,p149,p150,p151);
HA ha22(p120,p151,p152,p153);
FA fa54(p153,p122,p124,p154,p155);
FA fa55(ip_0_13,ip_1_12,ip_2_11,p156,p157);
FA fa56(ip_3_10,ip_4_9,ip_5_8,p158,p159);
FA fa57(ip_6_7,ip_7_6,ip_8_5,p160,p161);
HA ha23(ip_9_4,ip_10_3,p162,p163);
FA fa58(ip_11_2,ip_12_1,ip_13_0,p164,p165);
FA fa59(p126,p132,p163,p166,p167);
FA fa60(p157,p159,p161,p168,p169);
FA fa61(p165,p128,p130,p170,p171);
HA ha24(p134,p167,p172,p173);
FA fa62(p136,p140,p169,p174,p175);
FA fa63(p173,p138,p171,p176,p177);
FA fa64(p142,p146,p175,p178,p179);
FA fa65(p144,p177,p179,p180,p181);
HA ha25(p148,p181,p182,p183);
FA fa66(p150,p152,p183,p184,p185);
HA ha26(ip_0_14,ip_1_13,p186,p187);
FA fa67(ip_2_12,ip_3_11,ip_4_10,p188,p189);
FA fa68(ip_5_9,ip_6_8,ip_7_7,p190,p191);
FA fa69(ip_8_6,ip_9_5,ip_10_4,p192,p193);
FA fa70(ip_11_3,ip_12_2,ip_13_1,p194,p195);
FA fa71(ip_14_0,p162,p187,p196,p197);
FA fa72(p189,p191,p193,p198,p199);
FA fa73(p195,p156,p158,p200,p201);
FA fa74(p160,p164,p197,p202,p203);
FA fa75(p166,p172,p199,p204,p205);
FA fa76(p168,p201,p203,p206,p207);
FA fa77(p170,p205,p174,p208,p209);
FA fa78(p207,p176,p209,p210,p211);
FA fa79(p178,p180,p182,p212,p213);
FA fa80(p211,p213,p184,p214,p215);
FA fa81(ip_0_15,ip_1_14,ip_2_13,p216,p217);
FA fa82(ip_3_12,ip_4_11,ip_5_10,p218,p219);
FA fa83(ip_6_9,ip_7_8,ip_8_7,p220,p221);
FA fa84(ip_9_6,ip_10_5,ip_11_4,p222,p223);
FA fa85(ip_12_3,ip_13_2,ip_14_1,p224,p225);
HA ha27(ip_15_0,p186,p226,p227);
FA fa86(p217,p219,p221,p228,p229);
FA fa87(p223,p225,p227,p230,p231);
FA fa88(p188,p190,p192,p232,p233);
HA ha28(p194,p196,p234,p235);
FA fa89(p229,p231,p198,p236,p237);
FA fa90(p233,p235,p200,p238,p239);
FA fa91(p202,p237,p204,p240,p241);
FA fa92(p239,p206,p241,p242,p243);
HA ha29(p208,p243,p244,p245);
FA fa93(p210,p245,p212,p246,p247);
FA fa94(ip_0_16,ip_1_15,ip_2_14,p248,p249);
FA fa95(ip_3_13,ip_4_12,ip_5_11,p250,p251);
FA fa96(ip_6_10,ip_7_9,ip_8_8,p252,p253);
FA fa97(ip_9_7,ip_10_6,ip_11_5,p254,p255);
FA fa98(ip_12_4,ip_13_3,ip_14_2,p256,p257);
FA fa99(ip_15_1,ip_16_0,p226,p258,p259);
HA ha30(p249,p251,p260,p261);
HA ha31(p253,p255,p262,p263);
FA fa100(p257,p216,p218,p264,p265);
FA fa101(p220,p222,p224,p266,p267);
FA fa102(p259,p261,p263,p268,p269);
HA ha32(p228,p230,p270,p271);
FA fa103(p234,p265,p267,p272,p273);
FA fa104(p269,p232,p271,p274,p275);
FA fa105(p236,p273,p238,p276,p277);
FA fa106(p275,p240,p277,p278,p279);
FA fa107(p242,p244,p279,p280,p281);
FA fa108(ip_0_17,ip_1_16,ip_2_15,p282,p283);
FA fa109(ip_3_14,ip_4_13,ip_5_12,p284,p285);
FA fa110(ip_6_11,ip_7_10,ip_8_9,p286,p287);
FA fa111(ip_9_8,ip_10_7,ip_11_6,p288,p289);
FA fa112(ip_12_5,ip_13_4,ip_14_3,p290,p291);
FA fa113(ip_15_2,ip_16_1,ip_17_0,p292,p293);
FA fa114(p283,p285,p287,p294,p295);
FA fa115(p289,p291,p293,p296,p297);
FA fa116(p248,p250,p252,p298,p299);
FA fa117(p254,p256,p260,p300,p301);
FA fa118(p262,p258,p295,p302,p303);
HA ha33(p297,p299,p304,p305);
HA ha34(p301,p264,p306,p307);
HA ha35(p266,p268,p308,p309);
FA fa119(p270,p303,p305,p310,p311);
HA ha36(p307,p309,p312,p313);
HA ha37(p272,p311,p314,p315);
FA fa120(p313,p274,p315,p316,p317);
FA fa121(p276,p317,p278,p318,p319);
FA fa122(ip_0_18,ip_1_17,ip_2_16,p320,p321);
FA fa123(ip_3_15,ip_4_14,ip_5_13,p322,p323);
FA fa124(ip_6_12,ip_7_11,ip_8_10,p324,p325);
FA fa125(ip_9_9,ip_10_8,ip_11_7,p326,p327);
HA ha38(ip_12_6,ip_13_5,p328,p329);
FA fa126(ip_14_4,ip_15_3,ip_16_2,p330,p331);
FA fa127(ip_17_1,ip_18_0,p329,p332,p333);
HA ha39(p321,p323,p334,p335);
FA fa128(p325,p327,p331,p336,p337);
FA fa129(p333,p282,p284,p338,p339);
FA fa130(p286,p288,p290,p340,p341);
HA ha40(p292,p335,p342,p343);
HA ha41(p337,p343,p344,p345);
FA fa131(p294,p296,p339,p346,p347);
FA fa132(p341,p345,p298,p348,p349);
HA ha42(p300,p304,p350,p351);
FA fa133(p302,p306,p308,p352,p353);
FA fa134(p347,p349,p351,p354,p355);
FA fa135(p312,p310,p314,p356,p357);
FA fa136(p353,p355,p357,p358,p359);
FA fa137(p316,p359,p318,p360,p361);
FA fa138(ip_0_19,ip_1_18,ip_2_17,p362,p363);
FA fa139(ip_3_16,ip_4_15,ip_5_14,p364,p365);
FA fa140(ip_6_13,ip_7_12,ip_8_11,p366,p367);
FA fa141(ip_9_10,ip_10_9,ip_11_8,p368,p369);
FA fa142(ip_12_7,ip_13_6,ip_14_5,p370,p371);
FA fa143(ip_15_4,ip_16_3,ip_17_2,p372,p373);
FA fa144(ip_18_1,ip_19_0,p328,p374,p375);
FA fa145(p363,p365,p367,p376,p377);
FA fa146(p369,p371,p373,p378,p379);
FA fa147(p375,p320,p322,p380,p381);
HA ha43(p324,p326,p382,p383);
FA fa148(p330,p332,p334,p384,p385);
FA fa149(p342,p377,p379,p386,p387);
FA fa150(p383,p336,p344,p388,p389);
FA fa151(p381,p385,p338,p390,p391);
FA fa152(p340,p387,p350,p392,p393);
FA fa153(p389,p391,p346,p394,p395);
FA fa154(p348,p393,p395,p396,p397);
FA fa155(p352,p354,p397,p398,p399);
FA fa156(p356,p399,p358,p400,p401);
FA fa157(ip_0_20,ip_1_19,ip_2_18,p402,p403);
FA fa158(ip_3_17,ip_4_16,ip_5_15,p404,p405);
FA fa159(ip_6_14,ip_7_13,ip_8_12,p406,p407);
HA ha44(ip_9_11,ip_10_10,p408,p409);
FA fa160(ip_11_9,ip_12_8,ip_13_7,p410,p411);
FA fa161(ip_14_6,ip_15_5,ip_16_4,p412,p413);
FA fa162(ip_17_3,ip_18_2,ip_19_1,p414,p415);
FA fa163(ip_20_0,p409,p403,p416,p417);
HA ha45(p405,p407,p418,p419);
FA fa164(p411,p413,p415,p420,p421);
FA fa165(p362,p364,p366,p422,p423);
HA ha46(p368,p370,p424,p425);
FA fa166(p372,p374,p417,p426,p427);
FA fa167(p419,p382,p421,p428,p429);
FA fa168(p425,p376,p378,p430,p431);
FA fa169(p423,p427,p380,p432,p433);
FA fa170(p384,p429,p386,p434,p435);
FA fa171(p431,p433,p388,p436,p437);
HA ha47(p390,p435,p438,p439);
HA ha48(p392,p437,p440,p441);
HA ha49(p439,p394,p442,p443);
HA ha50(p441,p396,p444,p445);
FA fa172(p443,p445,p398,p446,p447);
FA fa173(ip_0_21,ip_1_20,ip_2_19,p448,p449);
HA ha51(ip_3_18,ip_4_17,p450,p451);
FA fa174(ip_5_16,ip_6_15,ip_7_14,p452,p453);
FA fa175(ip_8_13,ip_9_12,ip_10_11,p454,p455);
FA fa176(ip_11_10,ip_12_9,ip_13_8,p456,p457);
FA fa177(ip_14_7,ip_15_6,ip_16_5,p458,p459);
FA fa178(ip_17_4,ip_18_3,ip_19_2,p460,p461);
HA ha52(ip_20_1,ip_21_0,p462,p463);
FA fa179(p408,p451,p463,p464,p465);
FA fa180(p449,p453,p455,p466,p467);
HA ha53(p457,p459,p468,p469);
FA fa181(p461,p402,p404,p470,p471);
FA fa182(p406,p410,p412,p472,p473);
FA fa183(p414,p418,p465,p474,p475);
FA fa184(p469,p416,p424,p476,p477);
FA fa185(p467,p420,p471,p478,p479);
FA fa186(p473,p475,p422,p480,p481);
HA ha54(p426,p477,p482,p483);
HA ha55(p428,p479,p484,p485);
FA fa187(p481,p483,p430,p486,p487);
FA fa188(p432,p485,p434,p488,p489);
FA fa189(p438,p487,p436,p490,p491);
FA fa190(p440,p489,p442,p492,p493);
HA ha56(p491,p444,p494,p495);
FA fa191(p493,p495,p446,p496,p497);
FA fa192(ip_0_22,ip_1_21,ip_2_20,p498,p499);
FA fa193(ip_3_19,ip_4_18,ip_5_17,p500,p501);
HA ha57(ip_6_16,ip_7_15,p502,p503);
FA fa194(ip_8_14,ip_9_13,ip_10_12,p504,p505);
HA ha58(ip_11_11,ip_12_10,p506,p507);
HA ha59(ip_13_9,ip_14_8,p508,p509);
FA fa195(ip_15_7,ip_16_6,ip_17_5,p510,p511);
FA fa196(ip_18_4,ip_19_3,ip_20_2,p512,p513);
HA ha60(ip_21_1,ip_22_0,p514,p515);
FA fa197(p450,p462,p503,p516,p517);
FA fa198(p507,p509,p515,p518,p519);
FA fa199(p499,p501,p505,p520,p521);
FA fa200(p511,p513,p448,p522,p523);
HA ha61(p452,p454,p524,p525);
FA fa201(p456,p458,p460,p526,p527);
FA fa202(p468,p517,p519,p528,p529);
FA fa203(p464,p521,p523,p530,p531);
FA fa204(p525,p466,p527,p532,p533);
FA fa205(p529,p470,p472,p534,p535);
FA fa206(p474,p531,p476,p536,p537);
FA fa207(p482,p533,p478,p538,p539);
HA ha62(p480,p484,p540,p541);
FA fa208(p535,p537,p539,p542,p543);
HA ha63(p541,p486,p544,p545);
HA ha64(p543,p488,p546,p547);
FA fa209(p545,p490,p547,p548,p549);
FA fa210(p492,p494,p549,p550,p551);
FA fa211(ip_0_23,ip_1_22,ip_2_21,p552,p553);
FA fa212(ip_3_20,ip_4_19,ip_5_18,p554,p555);
FA fa213(ip_6_17,ip_7_16,ip_8_15,p556,p557);
HA ha65(ip_9_14,ip_10_13,p558,p559);
FA fa214(ip_11_12,ip_12_11,ip_13_10,p560,p561);
FA fa215(ip_14_9,ip_15_8,ip_16_7,p562,p563);
FA fa216(ip_17_6,ip_18_5,ip_19_4,p564,p565);
FA fa217(ip_20_3,ip_21_2,ip_22_1,p566,p567);
FA fa218(ip_23_0,p502,p506,p568,p569);
HA ha66(p508,p514,p570,p571);
HA ha67(p559,p553,p572,p573);
FA fa219(p555,p557,p561,p574,p575);
FA fa220(p563,p565,p567,p576,p577);
HA ha68(p571,p498,p578,p579);
FA fa221(p500,p504,p510,p580,p581);
FA fa222(p512,p569,p573,p582,p583);
FA fa223(p516,p518,p524,p584,p585);
FA fa224(p575,p577,p579,p586,p587);
FA fa225(p520,p522,p581,p588,p589);
FA fa226(p583,p526,p528,p590,p591);
FA fa227(p585,p587,p530,p592,p593);
FA fa228(p589,p532,p591,p594,p595);
FA fa229(p593,p534,p536,p596,p597);
FA fa230(p540,p538,p595,p598,p599);
FA fa231(p542,p544,p597,p600,p601);
FA fa232(p546,p599,p601,p602,p603);
FA fa233(p603,p548,p550,p604,p605);
FA fa234(ip_0_24,ip_1_23,ip_2_22,p606,p607);
FA fa235(ip_3_21,ip_4_20,ip_5_19,p608,p609);
FA fa236(ip_6_18,ip_7_17,ip_8_16,p610,p611);
FA fa237(ip_9_15,ip_10_14,ip_11_13,p612,p613);
FA fa238(ip_12_12,ip_13_11,ip_14_10,p614,p615);
FA fa239(ip_15_9,ip_16_8,ip_17_7,p616,p617);
FA fa240(ip_18_6,ip_19_5,ip_20_4,p618,p619);
HA ha69(ip_21_3,ip_22_2,p620,p621);
FA fa241(ip_23_1,ip_24_0,p558,p622,p623);
HA ha70(p621,p570,p624,p625);
FA fa242(p607,p609,p611,p626,p627);
HA ha71(p613,p615,p628,p629);
FA fa243(p617,p619,p623,p630,p631);
FA fa244(p552,p554,p556,p632,p633);
FA fa245(p560,p562,p564,p634,p635);
HA ha72(p566,p572,p636,p637);
FA fa246(p625,p629,p568,p638,p639);
HA ha73(p578,p627,p640,p641);
FA fa247(p631,p637,p574,p642,p643);
FA fa248(p576,p633,p635,p644,p645);
FA fa249(p639,p641,p580,p646,p647);
FA fa250(p582,p643,p584,p648,p649);
FA fa251(p586,p645,p647,p650,p651);
FA fa252(p588,p649,p590,p652,p653);
FA fa253(p592,p651,p653,p654,p655);
HA ha74(p594,p655,p656,p657);
FA fa254(p596,p657,p598,p658,p659);
FA fa255(p600,p659,p602,p660,p661);
FA fa256(ip_0_25,ip_1_24,ip_2_23,p662,p663);
FA fa257(ip_3_22,ip_4_21,ip_5_20,p664,p665);
FA fa258(ip_6_19,ip_7_18,ip_8_17,p666,p667);
FA fa259(ip_9_16,ip_10_15,ip_11_14,p668,p669);
FA fa260(ip_12_13,ip_13_12,ip_14_11,p670,p671);
FA fa261(ip_15_10,ip_16_9,ip_17_8,p672,p673);
FA fa262(ip_18_7,ip_19_6,ip_20_5,p674,p675);
FA fa263(ip_21_4,ip_22_3,ip_23_2,p676,p677);
FA fa264(ip_24_1,ip_25_0,p620,p678,p679);
FA fa265(p663,p665,p667,p680,p681);
FA fa266(p669,p671,p673,p682,p683);
HA ha75(p675,p677,p684,p685);
FA fa267(p679,p606,p608,p686,p687);
FA fa268(p610,p612,p614,p688,p689);
FA fa269(p616,p618,p622,p690,p691);
FA fa270(p624,p628,p685,p692,p693);
FA fa271(p636,p681,p683,p694,p695);
FA fa272(p626,p630,p640,p696,p697);
FA fa273(p687,p689,p691,p698,p699);
FA fa274(p693,p632,p634,p700,p701);
FA fa275(p638,p695,p642,p702,p703);
FA fa276(p697,p699,p644,p704,p705);
FA fa277(p646,p701,p703,p706,p707);
HA ha76(p648,p705,p708,p709);
FA fa278(p650,p707,p709,p710,p711);
HA ha77(p652,p654,p712,p713);
HA ha78(p656,p711,p714,p715);
FA fa279(p713,p715,p658,p716,p717);
FA fa280(ip_0_26,ip_1_25,ip_2_24,p718,p719);
FA fa281(ip_3_23,ip_4_22,ip_5_21,p720,p721);
HA ha79(ip_6_20,ip_7_19,p722,p723);
FA fa282(ip_8_18,ip_9_17,ip_10_16,p724,p725);
FA fa283(ip_11_15,ip_12_14,ip_13_13,p726,p727);
FA fa284(ip_14_12,ip_15_11,ip_16_10,p728,p729);
FA fa285(ip_17_9,ip_18_8,ip_19_7,p730,p731);
FA fa286(ip_20_6,ip_21_5,ip_22_4,p732,p733);
FA fa287(ip_23_3,ip_24_2,ip_25_1,p734,p735);
FA fa288(ip_26_0,p723,p719,p736,p737);
FA fa289(p721,p725,p727,p738,p739);
FA fa290(p729,p731,p733,p740,p741);
FA fa291(p735,p662,p664,p742,p743);
FA fa292(p666,p668,p670,p744,p745);
FA fa293(p672,p674,p676,p746,p747);
FA fa294(p678,p684,p737,p748,p749);
FA fa295(p739,p741,p680,p750,p751);
FA fa296(p682,p743,p745,p752,p753);
HA ha80(p747,p749,p754,p755);
FA fa297(p686,p688,p690,p756,p757);
FA fa298(p692,p751,p755,p758,p759);
FA fa299(p694,p753,p696,p760,p761);
FA fa300(p698,p757,p759,p762,p763);
FA fa301(p700,p702,p761,p764,p765);
FA fa302(p704,p708,p763,p766,p767);
HA ha81(p706,p765,p768,p769);
FA fa303(p767,p769,p710,p770,p771);
FA fa304(p712,p714,p771,p772,p773);
FA fa305(ip_0_27,ip_1_26,ip_2_25,p774,p775);
FA fa306(ip_3_24,ip_4_23,ip_5_22,p776,p777);
FA fa307(ip_6_21,ip_7_20,ip_8_19,p778,p779);
FA fa308(ip_9_18,ip_10_17,ip_11_16,p780,p781);
FA fa309(ip_12_15,ip_13_14,ip_14_13,p782,p783);
FA fa310(ip_15_12,ip_16_11,ip_17_10,p784,p785);
FA fa311(ip_18_9,ip_19_8,ip_20_7,p786,p787);
FA fa312(ip_21_6,ip_22_5,ip_23_4,p788,p789);
FA fa313(ip_24_3,ip_25_2,ip_26_1,p790,p791);
FA fa314(ip_27_0,p722,p775,p792,p793);
FA fa315(p777,p779,p781,p794,p795);
FA fa316(p783,p785,p787,p796,p797);
FA fa317(p789,p791,p718,p798,p799);
HA ha82(p720,p724,p800,p801);
HA ha83(p726,p728,p802,p803);
HA ha84(p730,p732,p804,p805);
FA fa318(p734,p793,p736,p806,p807);
HA ha85(p795,p797,p808,p809);
FA fa319(p799,p801,p803,p810,p811);
FA fa320(p805,p738,p740,p812,p813);
HA ha86(p807,p809,p814,p815);
FA fa321(p742,p744,p746,p816,p817);
FA fa322(p748,p754,p811,p818,p819);
HA ha87(p815,p750,p820,p821);
FA fa323(p813,p752,p817,p822,p823);
FA fa324(p819,p821,p756,p824,p825);
FA fa325(p758,p760,p823,p826,p827);
FA fa326(p825,p762,p764,p828,p829);
FA fa327(p768,p827,p766,p830,p831);
HA ha88(p829,p831,p832,p833);
FA fa328(p770,p833,p772,p834,p835);
FA fa329(ip_0_28,ip_1_27,ip_2_26,p836,p837);
HA ha89(ip_3_25,ip_4_24,p838,p839);
FA fa330(ip_5_23,ip_6_22,ip_7_21,p840,p841);
FA fa331(ip_8_20,ip_9_19,ip_10_18,p842,p843);
FA fa332(ip_11_17,ip_12_16,ip_13_15,p844,p845);
HA ha90(ip_14_14,ip_15_13,p846,p847);
FA fa333(ip_16_12,ip_17_11,ip_18_10,p848,p849);
FA fa334(ip_19_9,ip_20_8,ip_21_7,p850,p851);
FA fa335(ip_22_6,ip_23_5,ip_24_4,p852,p853);
FA fa336(ip_25_3,ip_26_2,ip_27_1,p854,p855);
FA fa337(ip_28_0,p839,p847,p856,p857);
HA ha91(p837,p841,p858,p859);
FA fa338(p843,p845,p849,p860,p861);
FA fa339(p851,p853,p855,p862,p863);
FA fa340(p774,p776,p778,p864,p865);
FA fa341(p780,p782,p784,p866,p867);
FA fa342(p786,p788,p790,p868,p869);
HA ha92(p857,p859,p870,p871);
HA ha93(p792,p800,p872,p873);
FA fa343(p802,p804,p861,p874,p875);
FA fa344(p863,p871,p794,p876,p877);
FA fa345(p796,p798,p808,p878,p879);
FA fa346(p865,p867,p869,p880,p881);
FA fa347(p873,p806,p814,p882,p883);
FA fa348(p875,p877,p810,p884,p885);
HA ha94(p879,p881,p886,p887);
FA fa349(p812,p820,p883,p888,p889);
HA ha95(p885,p887,p890,p891);
FA fa350(p816,p818,p891,p892,p893);
FA fa351(p889,p822,p824,p894,p895);
HA ha96(p893,p826,p896,p897);
FA fa352(p895,p828,p897,p898,p899);
FA fa353(p830,p832,p899,p900,p901);
FA fa354(ip_0_29,ip_1_28,ip_2_27,p902,p903);
HA ha97(ip_3_26,ip_4_25,p904,p905);
HA ha98(ip_5_24,ip_6_23,p906,p907);
HA ha99(ip_7_22,ip_8_21,p908,p909);
FA fa355(ip_9_20,ip_10_19,ip_11_18,p910,p911);
HA ha100(ip_12_17,ip_13_16,p912,p913);
HA ha101(ip_14_15,ip_15_14,p914,p915);
FA fa356(ip_16_13,ip_17_12,ip_18_11,p916,p917);
FA fa357(ip_19_10,ip_20_9,ip_21_8,p918,p919);
FA fa358(ip_22_7,ip_23_6,ip_24_5,p920,p921);
FA fa359(ip_25_4,ip_26_3,ip_27_2,p922,p923);
FA fa360(ip_28_1,ip_29_0,p838,p924,p925);
FA fa361(p846,p905,p907,p926,p927);
HA ha102(p909,p913,p928,p929);
FA fa362(p915,p903,p911,p930,p931);
FA fa363(p917,p919,p921,p932,p933);
FA fa364(p923,p925,p929,p934,p935);
HA ha103(p836,p840,p936,p937);
FA fa365(p842,p844,p848,p938,p939);
FA fa366(p850,p852,p854,p940,p941);
FA fa367(p858,p927,p856,p942,p943);
FA fa368(p870,p931,p933,p944,p945);
FA fa369(p935,p937,p860,p946,p947);
FA fa370(p862,p872,p939,p948,p949);
FA fa371(p941,p943,p864,p950,p951);
FA fa372(p866,p868,p945,p952,p953);
FA fa373(p947,p874,p876,p954,p955);
FA fa374(p949,p951,p878,p956,p957);
FA fa375(p880,p886,p953,p958,p959);
FA fa376(p882,p884,p890,p960,p961);
FA fa377(p955,p957,p959,p962,p963);
FA fa378(p888,p961,p963,p964,p965);
HA ha104(p892,p965,p966,p967);
FA fa379(p894,p896,p967,p968,p969);
FA fa380(p969,p898,p900,p970,p971);
FA fa381(ip_0_30,ip_1_29,ip_2_28,p972,p973);
HA ha105(ip_3_27,ip_4_26,p974,p975);
HA ha106(ip_5_25,ip_6_24,p976,p977);
FA fa382(ip_7_23,ip_8_22,ip_9_21,p978,p979);
FA fa383(ip_10_20,ip_11_19,ip_12_18,p980,p981);
FA fa384(ip_13_17,ip_14_16,ip_15_15,p982,p983);
HA ha107(ip_16_14,ip_17_13,p984,p985);
HA ha108(ip_18_12,ip_19_11,p986,p987);
FA fa385(ip_20_10,ip_21_9,ip_22_8,p988,p989);
FA fa386(ip_23_7,ip_24_6,ip_25_5,p990,p991);
HA ha109(ip_26_4,ip_27_3,p992,p993);
FA fa387(ip_28_2,ip_29_1,ip_30_0,p994,p995);
FA fa388(p904,p906,p908,p996,p997);
FA fa389(p912,p914,p975,p998,p999);
HA ha110(p977,p985,p1000,p1001);
HA ha111(p987,p993,p1002,p1003);
FA fa390(p1001,p1003,p928,p1004,p1005);
FA fa391(p973,p979,p981,p1006,p1007);
FA fa392(p983,p989,p991,p1008,p1009);
FA fa393(p995,p902,p910,p1010,p1011);
FA fa394(p916,p918,p920,p1012,p1013);
FA fa395(p922,p924,p997,p1014,p1015);
HA ha112(p999,p1005,p1016,p1017);
FA fa396(p1007,p1009,p926,p1018,p1019);
FA fa397(p936,p1011,p1013,p1020,p1021);
FA fa398(p1015,p1017,p930,p1022,p1023);
FA fa399(p932,p934,p1019,p1024,p1025);
FA fa400(p938,p940,p942,p1026,p1027);
FA fa401(p1021,p1023,p1025,p1028,p1029);
FA fa402(p944,p946,p1027,p1030,p1031);
FA fa403(p948,p950,p1029,p1032,p1033);
FA fa404(p1031,p952,p1033,p1034,p1035);
FA fa405(p954,p956,p1035,p1036,p1037);
FA fa406(p958,p1037,p960,p1038,p1039);
HA ha113(p962,p1039,p1040,p1041);
FA fa407(p964,p966,p1041,p1042,p1043);
FA fa408(p1043,p968,p970,p1044,p1045);
FA fa409(ip_0_31,ip_1_30,ip_2_29,p1046,p1047);
HA ha114(ip_3_28,ip_4_27,p1048,p1049);
FA fa410(ip_5_26,ip_6_25,ip_7_24,p1050,p1051);
FA fa411(ip_8_23,ip_9_22,ip_10_21,p1052,p1053);
FA fa412(ip_11_20,ip_12_19,ip_13_18,p1054,p1055);
FA fa413(ip_14_17,ip_15_16,ip_16_15,p1056,p1057);
FA fa414(ip_17_14,ip_18_13,ip_19_12,p1058,p1059);
FA fa415(ip_20_11,ip_21_10,ip_22_9,p1060,p1061);
FA fa416(ip_23_8,ip_24_7,ip_25_6,p1062,p1063);
FA fa417(ip_26_5,ip_27_4,ip_28_3,p1064,p1065);
FA fa418(ip_29_2,ip_30_1,ip_31_0,p1066,p1067);
FA fa419(p1049,p974,p976,p1068,p1069);
FA fa420(p984,p986,p992,p1070,p1071);
FA fa421(p1000,p1002,p1047,p1072,p1073);
HA ha115(p1051,p1053,p1074,p1075);
FA fa422(p1055,p1057,p1059,p1076,p1077);
FA fa423(p1061,p1063,p1065,p1078,p1079);
HA ha116(p1067,p1069,p1080,p1081);
FA fa424(p1071,p1075,p972,p1082,p1083);
FA fa425(p978,p980,p982,p1084,p1085);
FA fa426(p988,p990,p994,p1086,p1087);
FA fa427(p1073,p1077,p1079,p1088,p1089);
FA fa428(p1081,p996,p998,p1090,p1091);
FA fa429(p1004,p1006,p1008,p1092,p1093);
FA fa430(p1016,p1083,p1085,p1094,p1095);
FA fa431(p1087,p1010,p1012,p1096,p1097);
FA fa432(p1014,p1089,p1091,p1098,p1099);
FA fa433(p1018,p1093,p1095,p1100,p1101);
FA fa434(p1020,p1022,p1024,p1102,p1103);
FA fa435(p1097,p1099,p1026,p1104,p1105);
FA fa436(p1101,p1028,p1030,p1106,p1107);
FA fa437(p1103,p1105,p1032,p1108,p1109);
HA ha117(p1034,p1107,p1110,p1111);
FA fa438(p1109,p1036,p1111,p1112,p1113);
FA fa439(p1038,p1040,p1113,p1114,p1115);
FA fa440(p1042,p1115,p1044,p1116,p1117);
FA fa441(ip_0_32,ip_1_31,ip_2_30,p1118,p1119);
FA fa442(ip_3_29,ip_4_28,ip_5_27,p1120,p1121);
HA ha118(ip_6_26,ip_7_25,p1122,p1123);
HA ha119(ip_8_24,ip_9_23,p1124,p1125);
FA fa443(ip_10_22,ip_11_21,ip_12_20,p1126,p1127);
HA ha120(ip_13_19,ip_14_18,p1128,p1129);
FA fa444(ip_15_17,ip_16_16,ip_17_15,p1130,p1131);
HA ha121(ip_18_14,ip_19_13,p1132,p1133);
FA fa445(ip_20_12,ip_21_11,ip_22_10,p1134,p1135);
FA fa446(ip_23_9,ip_24_8,ip_25_7,p1136,p1137);
FA fa447(ip_26_6,ip_27_5,ip_28_4,p1138,p1139);
FA fa448(ip_29_3,ip_30_2,ip_31_1,p1140,p1141);
FA fa449(ip_32_0,p1048,p1123,p1142,p1143);
FA fa450(p1125,p1129,p1133,p1144,p1145);
FA fa451(p1119,p1121,p1127,p1146,p1147);
FA fa452(p1131,p1135,p1137,p1148,p1149);
FA fa453(p1139,p1141,p1046,p1150,p1151);
FA fa454(p1050,p1052,p1054,p1152,p1153);
HA ha122(p1056,p1058,p1154,p1155);
FA fa455(p1060,p1062,p1064,p1156,p1157);
FA fa456(p1066,p1074,p1143,p1158,p1159);
HA ha123(p1145,p1068,p1160,p1161);
HA ha124(p1070,p1080,p1162,p1163);
FA fa457(p1147,p1149,p1151,p1164,p1165);
FA fa458(p1155,p1072,p1076,p1166,p1167);
FA fa459(p1078,p1153,p1157,p1168,p1169);
HA ha125(p1159,p1161,p1170,p1171);
FA fa460(p1163,p1082,p1084,p1172,p1173);
FA fa461(p1086,p1165,p1171,p1174,p1175);
FA fa462(p1088,p1090,p1167,p1176,p1177);
FA fa463(p1169,p1092,p1094,p1178,p1179);
FA fa464(p1173,p1175,p1096,p1180,p1181);
FA fa465(p1098,p1177,p1100,p1182,p1183);
FA fa466(p1179,p1181,p1102,p1184,p1185);
FA fa467(p1104,p1183,p1185,p1186,p1187);
HA ha126(p1106,p1108,p1188,p1189);
FA fa468(p1110,p1187,p1189,p1190,p1191);
FA fa469(p1191,p1112,p1114,p1192,p1193);
HA ha127(ip_0_33,ip_1_32,p1194,p1195);
FA fa470(ip_2_31,ip_3_30,ip_4_29,p1196,p1197);
FA fa471(ip_5_28,ip_6_27,ip_7_26,p1198,p1199);
FA fa472(ip_8_25,ip_9_24,ip_10_23,p1200,p1201);
FA fa473(ip_11_22,ip_12_21,ip_13_20,p1202,p1203);
HA ha128(ip_14_19,ip_15_18,p1204,p1205);
FA fa474(ip_16_17,ip_17_16,ip_18_15,p1206,p1207);
FA fa475(ip_19_14,ip_20_13,ip_21_12,p1208,p1209);
FA fa476(ip_22_11,ip_23_10,ip_24_9,p1210,p1211);
HA ha129(ip_25_8,ip_26_7,p1212,p1213);
FA fa477(ip_27_6,ip_28_5,ip_29_4,p1214,p1215);
FA fa478(ip_30_3,ip_31_2,ip_32_1,p1216,p1217);
FA fa479(ip_33_0,p1122,p1124,p1218,p1219);
FA fa480(p1128,p1132,p1195,p1220,p1221);
FA fa481(p1205,p1213,p1197,p1222,p1223);
FA fa482(p1199,p1201,p1203,p1224,p1225);
FA fa483(p1207,p1209,p1211,p1226,p1227);
FA fa484(p1215,p1217,p1118,p1228,p1229);
FA fa485(p1120,p1126,p1130,p1230,p1231);
FA fa486(p1134,p1136,p1138,p1232,p1233);
HA ha130(p1140,p1219,p1234,p1235);
FA fa487(p1221,p1223,p1142,p1236,p1237);
FA fa488(p1144,p1154,p1225,p1238,p1239);
FA fa489(p1227,p1229,p1235,p1240,p1241);
FA fa490(p1146,p1148,p1150,p1242,p1243);
HA ha131(p1160,p1162,p1244,p1245);
HA ha132(p1231,p1233,p1246,p1247);
FA fa491(p1237,p1152,p1156,p1248,p1249);
FA fa492(p1158,p1170,p1239,p1250,p1251);
FA fa493(p1241,p1245,p1247,p1252,p1253);
FA fa494(p1164,p1243,p1166,p1254,p1255);
HA ha133(p1168,p1249,p1256,p1257);
FA fa495(p1251,p1253,p1172,p1258,p1259);
FA fa496(p1174,p1255,p1257,p1260,p1261);
FA fa497(p1176,p1259,p1178,p1262,p1263);
HA ha134(p1180,p1261,p1264,p1265);
FA fa498(p1182,p1263,p1265,p1266,p1267);
FA fa499(p1184,p1186,p1188,p1268,p1269);
FA fa500(p1267,p1190,p1269,p1270,p1271);
FA fa501(ip_0_34,ip_1_33,ip_2_32,p1272,p1273);
FA fa502(ip_3_31,ip_4_30,ip_5_29,p1274,p1275);
FA fa503(ip_6_28,ip_7_27,ip_8_26,p1276,p1277);
HA ha135(ip_9_25,ip_10_24,p1278,p1279);
FA fa504(ip_11_23,ip_12_22,ip_13_21,p1280,p1281);
HA ha136(ip_14_20,ip_15_19,p1282,p1283);
FA fa505(ip_16_18,ip_17_17,ip_18_16,p1284,p1285);
HA ha137(ip_19_15,ip_20_14,p1286,p1287);
FA fa506(ip_21_13,ip_22_12,ip_23_11,p1288,p1289);
FA fa507(ip_24_10,ip_25_9,ip_26_8,p1290,p1291);
HA ha138(ip_27_7,ip_28_6,p1292,p1293);
FA fa508(ip_29_5,ip_30_4,ip_31_3,p1294,p1295);
FA fa509(ip_32_2,ip_33_1,ip_34_0,p1296,p1297);
FA fa510(p1194,p1204,p1212,p1298,p1299);
FA fa511(p1279,p1283,p1287,p1300,p1301);
FA fa512(p1293,p1273,p1275,p1302,p1303);
FA fa513(p1277,p1281,p1285,p1304,p1305);
FA fa514(p1289,p1291,p1295,p1306,p1307);
FA fa515(p1297,p1196,p1198,p1308,p1309);
HA ha139(p1200,p1202,p1310,p1311);
FA fa516(p1206,p1208,p1210,p1312,p1313);
FA fa517(p1214,p1216,p1299,p1314,p1315);
FA fa518(p1301,p1218,p1220,p1316,p1317);
FA fa519(p1222,p1234,p1303,p1318,p1319);
FA fa520(p1305,p1307,p1311,p1320,p1321);
FA fa521(p1224,p1226,p1228,p1322,p1323);
HA ha140(p1309,p1313,p1324,p1325);
FA fa522(p1315,p1230,p1232,p1326,p1327);
FA fa523(p1236,p1244,p1246,p1328,p1329);
FA fa524(p1317,p1319,p1321,p1330,p1331);
HA ha141(p1325,p1238,p1332,p1333);
FA fa525(p1240,p1323,p1242,p1334,p1335);
FA fa526(p1327,p1329,p1331,p1336,p1337);
FA fa527(p1333,p1248,p1250,p1338,p1339);
FA fa528(p1252,p1256,p1335,p1340,p1341);
FA fa529(p1254,p1337,p1258,p1342,p1343);
HA ha142(p1339,p1341,p1344,p1345);
HA ha143(p1260,p1264,p1346,p1347);
HA ha144(p1343,p1345,p1348,p1349);
FA fa530(p1262,p1347,p1349,p1350,p1351);
FA fa531(p1266,p1351,p1268,p1352,p1353);
FA fa532(ip_0_35,ip_1_34,ip_2_33,p1354,p1355);
FA fa533(ip_3_32,ip_4_31,ip_5_30,p1356,p1357);
HA ha145(ip_6_29,ip_7_28,p1358,p1359);
FA fa534(ip_8_27,ip_9_26,ip_10_25,p1360,p1361);
FA fa535(ip_11_24,ip_12_23,ip_13_22,p1362,p1363);
HA ha146(ip_14_21,ip_15_20,p1364,p1365);
FA fa536(ip_16_19,ip_17_18,ip_18_17,p1366,p1367);
FA fa537(ip_19_16,ip_20_15,ip_21_14,p1368,p1369);
FA fa538(ip_22_13,ip_23_12,ip_24_11,p1370,p1371);
FA fa539(ip_25_10,ip_26_9,ip_27_8,p1372,p1373);
FA fa540(ip_28_7,ip_29_6,ip_30_5,p1374,p1375);
FA fa541(ip_31_4,ip_32_3,ip_33_2,p1376,p1377);
FA fa542(ip_34_1,ip_35_0,p1278,p1378,p1379);
FA fa543(p1282,p1286,p1292,p1380,p1381);
FA fa544(p1359,p1365,p1355,p1382,p1383);
FA fa545(p1357,p1361,p1363,p1384,p1385);
FA fa546(p1367,p1369,p1371,p1386,p1387);
FA fa547(p1373,p1375,p1377,p1388,p1389);
HA ha147(p1379,p1272,p1390,p1391);
HA ha148(p1274,p1276,p1392,p1393);
FA fa548(p1280,p1284,p1288,p1394,p1395);
FA fa549(p1290,p1294,p1296,p1396,p1397);
FA fa550(p1381,p1383,p1298,p1398,p1399);
FA fa551(p1300,p1310,p1385,p1400,p1401);
FA fa552(p1387,p1389,p1391,p1402,p1403);
HA ha149(p1393,p1302,p1404,p1405);
FA fa553(p1304,p1306,p1395,p1406,p1407);
FA fa554(p1397,p1399,p1308,p1408,p1409);
FA fa555(p1312,p1314,p1324,p1410,p1411);
HA ha150(p1401,p1403,p1412,p1413);
FA fa556(p1405,p1316,p1318,p1414,p1415);
FA fa557(p1320,p1407,p1409,p1416,p1417);
FA fa558(p1413,p1322,p1332,p1418,p1419);
FA fa559(p1411,p1326,p1328,p1420,p1421);
FA fa560(p1330,p1415,p1417,p1422,p1423);
FA fa561(p1334,p1419,p1336,p1424,p1425);
FA fa562(p1421,p1423,p1338,p1426,p1427);
HA ha151(p1340,p1344,p1428,p1429);
HA ha152(p1425,p1342,p1430,p1431);
FA fa563(p1346,p1348,p1427,p1432,p1433);
HA ha153(p1429,p1431,p1434,p1435);
FA fa564(p1433,p1435,p1350,p1436,p1437);
FA fa565(ip_0_36,ip_1_35,ip_2_34,p1438,p1439);
FA fa566(ip_3_33,ip_4_32,ip_5_31,p1440,p1441);
FA fa567(ip_6_30,ip_7_29,ip_8_28,p1442,p1443);
FA fa568(ip_9_27,ip_10_26,ip_11_25,p1444,p1445);
FA fa569(ip_12_24,ip_13_23,ip_14_22,p1446,p1447);
FA fa570(ip_15_21,ip_16_20,ip_17_19,p1448,p1449);
FA fa571(ip_18_18,ip_19_17,ip_20_16,p1450,p1451);
FA fa572(ip_21_15,ip_22_14,ip_23_13,p1452,p1453);
FA fa573(ip_24_12,ip_25_11,ip_26_10,p1454,p1455);
FA fa574(ip_27_9,ip_28_8,ip_29_7,p1456,p1457);
FA fa575(ip_30_6,ip_31_5,ip_32_4,p1458,p1459);
FA fa576(ip_33_3,ip_34_2,ip_35_1,p1460,p1461);
FA fa577(ip_36_0,p1358,p1364,p1462,p1463);
FA fa578(p1439,p1441,p1443,p1464,p1465);
FA fa579(p1445,p1447,p1449,p1466,p1467);
HA ha154(p1451,p1453,p1468,p1469);
FA fa580(p1455,p1457,p1459,p1470,p1471);
FA fa581(p1461,p1354,p1356,p1472,p1473);
HA ha155(p1360,p1362,p1474,p1475);
HA ha156(p1366,p1368,p1476,p1477);
FA fa582(p1370,p1372,p1374,p1478,p1479);
HA ha157(p1376,p1378,p1480,p1481);
HA ha158(p1463,p1469,p1482,p1483);
FA fa583(p1380,p1382,p1390,p1484,p1485);
FA fa584(p1392,p1465,p1467,p1486,p1487);
FA fa585(p1471,p1475,p1477,p1488,p1489);
HA ha159(p1481,p1483,p1490,p1491);
FA fa586(p1384,p1386,p1388,p1492,p1493);
FA fa587(p1473,p1479,p1491,p1494,p1495);
HA ha160(p1394,p1396,p1496,p1497);
FA fa588(p1398,p1404,p1485,p1498,p1499);
HA ha161(p1487,p1489,p1500,p1501);
HA ha162(p1400,p1402,p1502,p1503);
FA fa589(p1412,p1493,p1495,p1504,p1505);
HA ha163(p1497,p1501,p1506,p1507);
FA fa590(p1406,p1408,p1499,p1508,p1509);
FA fa591(p1503,p1507,p1410,p1510,p1511);
FA fa592(p1505,p1414,p1416,p1512,p1513);
FA fa593(p1509,p1511,p1418,p1514,p1515);
FA fa594(p1420,p1422,p1513,p1516,p1517);
FA fa595(p1515,p1424,p1428,p1518,p1519);
FA fa596(p1426,p1430,p1517,p1520,p1521);
HA ha164(p1434,p1519,p1522,p1523);
FA fa597(p1432,p1521,p1523,p1524,p1525);
FA fa598(ip_0_37,ip_1_36,ip_2_35,p1526,p1527);
FA fa599(ip_3_34,ip_4_33,ip_5_32,p1528,p1529);
FA fa600(ip_6_31,ip_7_30,ip_8_29,p1530,p1531);
FA fa601(ip_9_28,ip_10_27,ip_11_26,p1532,p1533);
FA fa602(ip_12_25,ip_13_24,ip_14_23,p1534,p1535);
FA fa603(ip_15_22,ip_16_21,ip_17_20,p1536,p1537);
HA ha165(ip_18_19,ip_19_18,p1538,p1539);
FA fa604(ip_20_17,ip_21_16,ip_22_15,p1540,p1541);
FA fa605(ip_23_14,ip_24_13,ip_25_12,p1542,p1543);
FA fa606(ip_26_11,ip_27_10,ip_28_9,p1544,p1545);
FA fa607(ip_29_8,ip_30_7,ip_31_6,p1546,p1547);
FA fa608(ip_32_5,ip_33_4,ip_34_3,p1548,p1549);
HA ha166(ip_35_2,ip_36_1,p1550,p1551);
FA fa609(ip_37_0,p1539,p1551,p1552,p1553);
FA fa610(p1527,p1529,p1531,p1554,p1555);
HA ha167(p1533,p1535,p1556,p1557);
FA fa611(p1537,p1541,p1543,p1558,p1559);
FA fa612(p1545,p1547,p1549,p1560,p1561);
HA ha168(p1438,p1440,p1562,p1563);
HA ha169(p1442,p1444,p1564,p1565);
FA fa613(p1446,p1448,p1450,p1566,p1567);
FA fa614(p1452,p1454,p1456,p1568,p1569);
FA fa615(p1458,p1460,p1468,p1570,p1571);
HA ha170(p1553,p1557,p1572,p1573);
FA fa616(p1462,p1474,p1476,p1574,p1575);
FA fa617(p1480,p1482,p1555,p1576,p1577);
FA fa618(p1559,p1561,p1563,p1578,p1579);
FA fa619(p1565,p1573,p1464,p1580,p1581);
HA ha171(p1466,p1470,p1582,p1583);
FA fa620(p1490,p1567,p1569,p1584,p1585);
FA fa621(p1571,p1472,p1478,p1586,p1587);
FA fa622(p1575,p1577,p1579,p1588,p1589);
FA fa623(p1581,p1583,p1484,p1590,p1591);
FA fa624(p1486,p1488,p1496,p1592,p1593);
FA fa625(p1500,p1585,p1492,p1594,p1595);
FA fa626(p1494,p1502,p1506,p1596,p1597);
FA fa627(p1587,p1589,p1591,p1598,p1599);
FA fa628(p1498,p1593,p1595,p1600,p1601);
FA fa629(p1504,p1597,p1599,p1602,p1603);
FA fa630(p1508,p1510,p1601,p1604,p1605);
FA fa631(p1603,p1512,p1514,p1606,p1607);
FA fa632(p1605,p1516,p1607,p1608,p1609);
HA ha172(p1518,p1522,p1610,p1611);
HA ha173(p1520,p1609,p1612,p1613);
FA fa633(p1611,p1613,p1524,p1614,p1615);
FA fa634(ip_0_38,ip_1_37,ip_2_36,p1616,p1617);
FA fa635(ip_3_35,ip_4_34,ip_5_33,p1618,p1619);
FA fa636(ip_6_32,ip_7_31,ip_8_30,p1620,p1621);
FA fa637(ip_9_29,ip_10_28,ip_11_27,p1622,p1623);
FA fa638(ip_12_26,ip_13_25,ip_14_24,p1624,p1625);
FA fa639(ip_15_23,ip_16_22,ip_17_21,p1626,p1627);
FA fa640(ip_18_20,ip_19_19,ip_20_18,p1628,p1629);
FA fa641(ip_21_17,ip_22_16,ip_23_15,p1630,p1631);
FA fa642(ip_24_14,ip_25_13,ip_26_12,p1632,p1633);
FA fa643(ip_27_11,ip_28_10,ip_29_9,p1634,p1635);
FA fa644(ip_30_8,ip_31_7,ip_32_6,p1636,p1637);
FA fa645(ip_33_5,ip_34_4,ip_35_3,p1638,p1639);
HA ha174(ip_36_2,ip_37_1,p1640,p1641);
FA fa646(ip_38_0,p1538,p1550,p1642,p1643);
HA ha175(p1641,p1617,p1644,p1645);
FA fa647(p1619,p1621,p1623,p1646,p1647);
FA fa648(p1625,p1627,p1629,p1648,p1649);
FA fa649(p1631,p1633,p1635,p1650,p1651);
FA fa650(p1637,p1639,p1526,p1652,p1653);
FA fa651(p1528,p1530,p1532,p1654,p1655);
FA fa652(p1534,p1536,p1540,p1656,p1657);
HA ha176(p1542,p1544,p1658,p1659);
FA fa653(p1546,p1548,p1556,p1660,p1661);
FA fa654(p1643,p1645,p1552,p1662,p1663);
FA fa655(p1562,p1564,p1572,p1664,p1665);
FA fa656(p1647,p1649,p1651,p1666,p1667);
FA fa657(p1653,p1659,p1554,p1668,p1669);
FA fa658(p1558,p1560,p1655,p1670,p1671);
FA fa659(p1657,p1661,p1663,p1672,p1673);
HA ha177(p1566,p1568,p1674,p1675);
FA fa660(p1570,p1582,p1665,p1676,p1677);
FA fa661(p1667,p1669,p1574,p1678,p1679);
FA fa662(p1576,p1578,p1580,p1680,p1681);
FA fa663(p1671,p1673,p1675,p1682,p1683);
HA ha178(p1584,p1677,p1684,p1685);
FA fa664(p1679,p1586,p1588,p1686,p1687);
FA fa665(p1590,p1681,p1683,p1688,p1689);
FA fa666(p1685,p1592,p1594,p1690,p1691);
FA fa667(p1596,p1598,p1687,p1692,p1693);
FA fa668(p1689,p1600,p1691,p1694,p1695);
HA ha179(p1602,p1693,p1696,p1697);
FA fa669(p1604,p1695,p1697,p1698,p1699);
FA fa670(p1606,p1699,p1610,p1700,p1701);
FA fa671(p1608,p1612,p1701,p1702,p1703);
FA fa672(ip_0_39,ip_1_38,ip_2_37,p1704,p1705);
FA fa673(ip_3_36,ip_4_35,ip_5_34,p1706,p1707);
FA fa674(ip_6_33,ip_7_32,ip_8_31,p1708,p1709);
FA fa675(ip_9_30,ip_10_29,ip_11_28,p1710,p1711);
FA fa676(ip_12_27,ip_13_26,ip_14_25,p1712,p1713);
FA fa677(ip_15_24,ip_16_23,ip_17_22,p1714,p1715);
FA fa678(ip_18_21,ip_19_20,ip_20_19,p1716,p1717);
HA ha180(ip_21_18,ip_22_17,p1718,p1719);
FA fa679(ip_23_16,ip_24_15,ip_25_14,p1720,p1721);
FA fa680(ip_26_13,ip_27_12,ip_28_11,p1722,p1723);
FA fa681(ip_29_10,ip_30_9,ip_31_8,p1724,p1725);
FA fa682(ip_32_7,ip_33_6,ip_34_5,p1726,p1727);
FA fa683(ip_35_4,ip_36_3,ip_37_2,p1728,p1729);
FA fa684(ip_38_1,ip_39_0,p1640,p1730,p1731);
FA fa685(p1719,p1705,p1707,p1732,p1733);
FA fa686(p1709,p1711,p1713,p1734,p1735);
FA fa687(p1715,p1717,p1721,p1736,p1737);
FA fa688(p1723,p1725,p1727,p1738,p1739);
FA fa689(p1729,p1731,p1616,p1740,p1741);
FA fa690(p1618,p1620,p1622,p1742,p1743);
FA fa691(p1624,p1626,p1628,p1744,p1745);
FA fa692(p1630,p1632,p1634,p1746,p1747);
FA fa693(p1636,p1638,p1644,p1748,p1749);
HA ha181(p1642,p1658,p1750,p1751);
FA fa694(p1733,p1735,p1737,p1752,p1753);
FA fa695(p1739,p1741,p1646,p1754,p1755);
HA ha182(p1648,p1650,p1756,p1757);
FA fa696(p1652,p1743,p1745,p1758,p1759);
FA fa697(p1747,p1749,p1751,p1760,p1761);
FA fa698(p1654,p1656,p1660,p1762,p1763);
FA fa699(p1662,p1753,p1755,p1764,p1765);
FA fa700(p1757,p1664,p1666,p1766,p1767);
FA fa701(p1668,p1674,p1759,p1768,p1769);
FA fa702(p1761,p1670,p1672,p1770,p1771);
FA fa703(p1763,p1765,p1676,p1772,p1773);
HA ha183(p1678,p1684,p1774,p1775);
HA ha184(p1767,p1769,p1776,p1777);
FA fa704(p1680,p1682,p1771,p1778,p1779);
FA fa705(p1773,p1775,p1777,p1780,p1781);
FA fa706(p1686,p1688,p1779,p1782,p1783);
FA fa707(p1781,p1690,p1692,p1784,p1785);
FA fa708(p1696,p1783,p1694,p1786,p1787);
FA fa709(p1785,p1787,p1698,p1788,p1789);
FA fa710(p1789,p1700,p1702,p1790,p1791);
FA fa711(ip_0_40,ip_1_39,ip_2_38,p1792,p1793);
FA fa712(ip_3_37,ip_4_36,ip_5_35,p1794,p1795);
FA fa713(ip_6_34,ip_7_33,ip_8_32,p1796,p1797);
FA fa714(ip_9_31,ip_10_30,ip_11_29,p1798,p1799);
FA fa715(ip_12_28,ip_13_27,ip_14_26,p1800,p1801);
FA fa716(ip_15_25,ip_16_24,ip_17_23,p1802,p1803);
FA fa717(ip_18_22,ip_19_21,ip_20_20,p1804,p1805);
FA fa718(ip_21_19,ip_22_18,ip_23_17,p1806,p1807);
FA fa719(ip_24_16,ip_25_15,ip_26_14,p1808,p1809);
FA fa720(ip_27_13,ip_28_12,ip_29_11,p1810,p1811);
FA fa721(ip_30_10,ip_31_9,ip_32_8,p1812,p1813);
FA fa722(ip_33_7,ip_34_6,ip_35_5,p1814,p1815);
FA fa723(ip_36_4,ip_37_3,ip_38_2,p1816,p1817);
FA fa724(ip_39_1,ip_40_0,p1718,p1818,p1819);
FA fa725(p1793,p1795,p1797,p1820,p1821);
FA fa726(p1799,p1801,p1803,p1822,p1823);
FA fa727(p1805,p1807,p1809,p1824,p1825);
FA fa728(p1811,p1813,p1815,p1826,p1827);
FA fa729(p1817,p1819,p1704,p1828,p1829);
HA ha185(p1706,p1708,p1830,p1831);
HA ha186(p1710,p1712,p1832,p1833);
FA fa730(p1714,p1716,p1720,p1834,p1835);
FA fa731(p1722,p1724,p1726,p1836,p1837);
FA fa732(p1728,p1730,p1821,p1838,p1839);
FA fa733(p1823,p1825,p1827,p1840,p1841);
FA fa734(p1829,p1831,p1833,p1842,p1843);
FA fa735(p1732,p1734,p1736,p1844,p1845);
FA fa736(p1738,p1740,p1750,p1846,p1847);
FA fa737(p1835,p1837,p1839,p1848,p1849);
FA fa738(p1742,p1744,p1746,p1850,p1851);
FA fa739(p1748,p1756,p1841,p1852,p1853);
FA fa740(p1843,p1752,p1754,p1854,p1855);
FA fa741(p1845,p1847,p1849,p1856,p1857);
FA fa742(p1758,p1760,p1851,p1858,p1859);
FA fa743(p1853,p1762,p1764,p1860,p1861);
FA fa744(p1855,p1857,p1766,p1862,p1863);
FA fa745(p1768,p1774,p1776,p1864,p1865);
FA fa746(p1859,p1770,p1772,p1866,p1867);
FA fa747(p1861,p1863,p1865,p1868,p1869);
FA fa748(p1778,p1780,p1867,p1870,p1871);
HA ha187(p1869,p1782,p1872,p1873);
FA fa749(p1871,p1784,p1873,p1874,p1875);
FA fa750(p1786,p1875,p1788,p1876,p1877);
FA fa751(ip_0_41,ip_1_40,ip_2_39,p1878,p1879);
HA ha188(ip_3_38,ip_4_37,p1880,p1881);
FA fa752(ip_5_36,ip_6_35,ip_7_34,p1882,p1883);
FA fa753(ip_8_33,ip_9_32,ip_10_31,p1884,p1885);
FA fa754(ip_11_30,ip_12_29,ip_13_28,p1886,p1887);
FA fa755(ip_14_27,ip_15_26,ip_16_25,p1888,p1889);
FA fa756(ip_17_24,ip_18_23,ip_19_22,p1890,p1891);
FA fa757(ip_20_21,ip_21_20,ip_22_19,p1892,p1893);
FA fa758(ip_23_18,ip_24_17,ip_25_16,p1894,p1895);
FA fa759(ip_26_15,ip_27_14,ip_28_13,p1896,p1897);
HA ha189(ip_29_12,ip_30_11,p1898,p1899);
FA fa760(ip_31_10,ip_32_9,ip_33_8,p1900,p1901);
FA fa761(ip_34_7,ip_35_6,ip_36_5,p1902,p1903);
FA fa762(ip_37_4,ip_38_3,ip_39_2,p1904,p1905);
FA fa763(ip_40_1,ip_41_0,p1881,p1906,p1907);
FA fa764(p1899,p1879,p1883,p1908,p1909);
HA ha190(p1885,p1887,p1910,p1911);
HA ha191(p1889,p1891,p1912,p1913);
FA fa765(p1893,p1895,p1897,p1914,p1915);
FA fa766(p1901,p1903,p1905,p1916,p1917);
FA fa767(p1907,p1792,p1794,p1918,p1919);
FA fa768(p1796,p1798,p1800,p1920,p1921);
HA ha192(p1802,p1804,p1922,p1923);
FA fa769(p1806,p1808,p1810,p1924,p1925);
FA fa770(p1812,p1814,p1816,p1926,p1927);
FA fa771(p1818,p1911,p1913,p1928,p1929);
FA fa772(p1830,p1832,p1909,p1930,p1931);
FA fa773(p1915,p1917,p1923,p1932,p1933);
HA ha193(p1820,p1822,p1934,p1935);
FA fa774(p1824,p1826,p1828,p1936,p1937);
HA ha194(p1919,p1921,p1938,p1939);
FA fa775(p1925,p1927,p1929,p1940,p1941);
FA fa776(p1834,p1836,p1838,p1942,p1943);
FA fa777(p1931,p1933,p1935,p1944,p1945);
FA fa778(p1939,p1840,p1842,p1946,p1947);
FA fa779(p1937,p1941,p1844,p1948,p1949);
HA ha195(p1846,p1848,p1950,p1951);
FA fa780(p1943,p1945,p1850,p1952,p1953);
FA fa781(p1852,p1947,p1949,p1954,p1955);
HA ha196(p1951,p1854,p1956,p1957);
FA fa782(p1856,p1953,p1858,p1958,p1959);
FA fa783(p1955,p1957,p1860,p1960,p1961);
HA ha197(p1862,p1959,p1962,p1963);
FA fa784(p1864,p1961,p1963,p1964,p1965);
FA fa785(p1866,p1868,p1965,p1966,p1967);
FA fa786(p1870,p1872,p1967,p1968,p1969);
HA ha198(p1969,p1874,p1970,p1971);
HA ha199(ip_0_42,ip_1_41,p1972,p1973);
FA fa787(ip_2_40,ip_3_39,ip_4_38,p1974,p1975);
FA fa788(ip_5_37,ip_6_36,ip_7_35,p1976,p1977);
FA fa789(ip_8_34,ip_9_33,ip_10_32,p1978,p1979);
FA fa790(ip_11_31,ip_12_30,ip_13_29,p1980,p1981);
FA fa791(ip_14_28,ip_15_27,ip_16_26,p1982,p1983);
FA fa792(ip_17_25,ip_18_24,ip_19_23,p1984,p1985);
FA fa793(ip_20_22,ip_21_21,ip_22_20,p1986,p1987);
FA fa794(ip_23_19,ip_24_18,ip_25_17,p1988,p1989);
FA fa795(ip_26_16,ip_27_15,ip_28_14,p1990,p1991);
FA fa796(ip_29_13,ip_30_12,ip_31_11,p1992,p1993);
HA ha200(ip_32_10,ip_33_9,p1994,p1995);
FA fa797(ip_34_8,ip_35_7,ip_36_6,p1996,p1997);
FA fa798(ip_37_5,ip_38_4,ip_39_3,p1998,p1999);
FA fa799(ip_40_2,ip_41_1,ip_42_0,p2000,p2001);
FA fa800(p1880,p1898,p1973,p2002,p2003);
FA fa801(p1995,p1975,p1977,p2004,p2005);
FA fa802(p1979,p1981,p1983,p2006,p2007);
HA ha201(p1985,p1987,p2008,p2009);
FA fa803(p1989,p1991,p1993,p2010,p2011);
FA fa804(p1997,p1999,p2001,p2012,p2013);
FA fa805(p1878,p1882,p1884,p2014,p2015);
FA fa806(p1886,p1888,p1890,p2016,p2017);
FA fa807(p1892,p1894,p1896,p2018,p2019);
HA ha202(p1900,p1902,p2020,p2021);
HA ha203(p1904,p1906,p2022,p2023);
FA fa808(p1910,p1912,p2003,p2024,p2025);
FA fa809(p2009,p1922,p2005,p2026,p2027);
FA fa810(p2007,p2011,p2013,p2028,p2029);
FA fa811(p2021,p2023,p1908,p2030,p2031);
FA fa812(p1914,p1916,p2015,p2032,p2033);
FA fa813(p2017,p2019,p2025,p2034,p2035);
FA fa814(p1918,p1920,p1924,p2036,p2037);
FA fa815(p1926,p1928,p1934,p2038,p2039);
FA fa816(p1938,p2027,p2029,p2040,p2041);
HA ha204(p2031,p1930,p2042,p2043);
FA fa817(p1932,p2033,p2035,p2044,p2045);
FA fa818(p1936,p1940,p2037,p2046,p2047);
HA ha205(p2039,p2041,p2048,p2049);
FA fa819(p2043,p1942,p1944,p2050,p2051);
FA fa820(p1950,p2045,p2049,p2052,p2053);
FA fa821(p1946,p1948,p2047,p2054,p2055);
FA fa822(p1952,p1956,p2051,p2056,p2057);
FA fa823(p2053,p1954,p2055,p2058,p2059);
FA fa824(p1958,p1962,p2057,p2060,p2061);
FA fa825(p1960,p2059,p2061,p2062,p2063);
HA ha206(p1964,p2063,p2064,p2065);
HA ha207(p1966,p2065,p2066,p2067);
FA fa826(p2067,p1968,p1970,p2068,p2069);
FA fa827(ip_0_43,ip_1_42,ip_2_41,p2070,p2071);
HA ha208(ip_3_40,ip_4_39,p2072,p2073);
FA fa828(ip_5_38,ip_6_37,ip_7_36,p2074,p2075);
FA fa829(ip_8_35,ip_9_34,ip_10_33,p2076,p2077);
HA ha209(ip_11_32,ip_12_31,p2078,p2079);
FA fa830(ip_13_30,ip_14_29,ip_15_28,p2080,p2081);
FA fa831(ip_16_27,ip_17_26,ip_18_25,p2082,p2083);
FA fa832(ip_19_24,ip_20_23,ip_21_22,p2084,p2085);
FA fa833(ip_22_21,ip_23_20,ip_24_19,p2086,p2087);
FA fa834(ip_25_18,ip_26_17,ip_27_16,p2088,p2089);
FA fa835(ip_28_15,ip_29_14,ip_30_13,p2090,p2091);
FA fa836(ip_31_12,ip_32_11,ip_33_10,p2092,p2093);
FA fa837(ip_34_9,ip_35_8,ip_36_7,p2094,p2095);
FA fa838(ip_37_6,ip_38_5,ip_39_4,p2096,p2097);
FA fa839(ip_40_3,ip_41_2,ip_42_1,p2098,p2099);
FA fa840(ip_43_0,p1972,p1994,p2100,p2101);
FA fa841(p2073,p2079,p2071,p2102,p2103);
HA ha210(p2075,p2077,p2104,p2105);
FA fa842(p2081,p2083,p2085,p2106,p2107);
FA fa843(p2087,p2089,p2091,p2108,p2109);
HA ha211(p2093,p2095,p2110,p2111);
FA fa844(p2097,p2099,p1974,p2112,p2113);
FA fa845(p1976,p1978,p1980,p2114,p2115);
FA fa846(p1982,p1984,p1986,p2116,p2117);
FA fa847(p1988,p1990,p1992,p2118,p2119);
FA fa848(p1996,p1998,p2000,p2120,p2121);
FA fa849(p2008,p2101,p2103,p2122,p2123);
FA fa850(p2105,p2111,p2002,p2124,p2125);
FA fa851(p2020,p2022,p2107,p2126,p2127);
FA fa852(p2109,p2113,p2004,p2128,p2129);
FA fa853(p2006,p2010,p2012,p2130,p2131);
FA fa854(p2115,p2117,p2119,p2132,p2133);
FA fa855(p2121,p2123,p2125,p2134,p2135);
HA ha212(p2014,p2016,p2136,p2137);
FA fa856(p2018,p2024,p2127,p2138,p2139);
FA fa857(p2129,p2026,p2028,p2140,p2141);
HA ha213(p2030,p2131,p2142,p2143);
FA fa858(p2133,p2135,p2137,p2144,p2145);
HA ha214(p2032,p2034,p2146,p2147);
FA fa859(p2042,p2139,p2143,p2148,p2149);
FA fa860(p2036,p2038,p2040,p2150,p2151);
FA fa861(p2048,p2141,p2145,p2152,p2153);
FA fa862(p2147,p2044,p2149,p2154,p2155);
HA ha215(p2046,p2151,p2156,p2157);
FA fa863(p2153,p2050,p2052,p2158,p2159);
FA fa864(p2155,p2157,p2054,p2160,p2161);
HA ha216(p2056,p2159,p2162,p2163);
FA fa865(p2161,p2058,p2163,p2164,p2165);
FA fa866(p2060,p2062,p2064,p2166,p2167);
FA fa867(p2165,p2066,p2167,p2168,p2169);
FA fa868(ip_0_44,ip_1_43,ip_2_42,p2170,p2171);
FA fa869(ip_3_41,ip_4_40,ip_5_39,p2172,p2173);
HA ha217(ip_6_38,ip_7_37,p2174,p2175);
FA fa870(ip_8_36,ip_9_35,ip_10_34,p2176,p2177);
FA fa871(ip_11_33,ip_12_32,ip_13_31,p2178,p2179);
FA fa872(ip_14_30,ip_15_29,ip_16_28,p2180,p2181);
FA fa873(ip_17_27,ip_18_26,ip_19_25,p2182,p2183);
FA fa874(ip_20_24,ip_21_23,ip_22_22,p2184,p2185);
HA ha218(ip_23_21,ip_24_20,p2186,p2187);
HA ha219(ip_25_19,ip_26_18,p2188,p2189);
FA fa875(ip_27_17,ip_28_16,ip_29_15,p2190,p2191);
HA ha220(ip_30_14,ip_31_13,p2192,p2193);
HA ha221(ip_32_12,ip_33_11,p2194,p2195);
FA fa876(ip_34_10,ip_35_9,ip_36_8,p2196,p2197);
FA fa877(ip_37_7,ip_38_6,ip_39_5,p2198,p2199);
FA fa878(ip_40_4,ip_41_3,ip_42_2,p2200,p2201);
FA fa879(ip_43_1,ip_44_0,p2072,p2202,p2203);
FA fa880(p2078,p2175,p2187,p2204,p2205);
FA fa881(p2189,p2193,p2195,p2206,p2207);
HA ha222(p2171,p2173,p2208,p2209);
FA fa882(p2177,p2179,p2181,p2210,p2211);
HA ha223(p2183,p2185,p2212,p2213);
FA fa883(p2191,p2197,p2199,p2214,p2215);
FA fa884(p2201,p2203,p2070,p2216,p2217);
FA fa885(p2074,p2076,p2080,p2218,p2219);
FA fa886(p2082,p2084,p2086,p2220,p2221);
FA fa887(p2088,p2090,p2092,p2222,p2223);
HA ha224(p2094,p2096,p2224,p2225);
FA fa888(p2098,p2104,p2110,p2226,p2227);
HA ha225(p2205,p2207,p2228,p2229);
FA fa889(p2209,p2213,p2100,p2230,p2231);
HA ha226(p2102,p2211,p2232,p2233);
FA fa890(p2215,p2217,p2225,p2234,p2235);
HA ha227(p2229,p2106,p2236,p2237);
FA fa891(p2108,p2112,p2219,p2238,p2239);
FA fa892(p2221,p2223,p2227,p2240,p2241);
FA fa893(p2231,p2233,p2114,p2242,p2243);
FA fa894(p2116,p2118,p2120,p2244,p2245);
FA fa895(p2122,p2124,p2235,p2246,p2247);
FA fa896(p2237,p2126,p2128,p2248,p2249);
FA fa897(p2136,p2239,p2241,p2250,p2251);
FA fa898(p2243,p2130,p2132,p2252,p2253);
FA fa899(p2134,p2142,p2245,p2254,p2255);
FA fa900(p2247,p2138,p2146,p2256,p2257);
FA fa901(p2249,p2251,p2140,p2258,p2259);
FA fa902(p2144,p2253,p2255,p2260,p2261);
FA fa903(p2148,p2257,p2259,p2262,p2263);
FA fa904(p2150,p2152,p2156,p2264,p2265);
FA fa905(p2261,p2154,p2263,p2266,p2267);
FA fa906(p2265,p2158,p2160,p2268,p2269);
FA fa907(p2162,p2267,p2269,p2270,p2271);
FA fa908(p2164,p2271,p2166,p2272,p2273);
FA fa909(ip_0_45,ip_1_44,ip_2_43,p2274,p2275);
FA fa910(ip_3_42,ip_4_41,ip_5_40,p2276,p2277);
FA fa911(ip_6_39,ip_7_38,ip_8_37,p2278,p2279);
FA fa912(ip_9_36,ip_10_35,ip_11_34,p2280,p2281);
HA ha228(ip_12_33,ip_13_32,p2282,p2283);
FA fa913(ip_14_31,ip_15_30,ip_16_29,p2284,p2285);
FA fa914(ip_17_28,ip_18_27,ip_19_26,p2286,p2287);
HA ha229(ip_20_25,ip_21_24,p2288,p2289);
FA fa915(ip_22_23,ip_23_22,ip_24_21,p2290,p2291);
FA fa916(ip_25_20,ip_26_19,ip_27_18,p2292,p2293);
FA fa917(ip_28_17,ip_29_16,ip_30_15,p2294,p2295);
FA fa918(ip_31_14,ip_32_13,ip_33_12,p2296,p2297);
FA fa919(ip_34_11,ip_35_10,ip_36_9,p2298,p2299);
FA fa920(ip_37_8,ip_38_7,ip_39_6,p2300,p2301);
HA ha230(ip_40_5,ip_41_4,p2302,p2303);
FA fa921(ip_42_3,ip_43_2,ip_44_1,p2304,p2305);
FA fa922(ip_45_0,p2174,p2186,p2306,p2307);
FA fa923(p2188,p2192,p2194,p2308,p2309);
FA fa924(p2283,p2289,p2303,p2310,p2311);
FA fa925(p2275,p2277,p2279,p2312,p2313);
FA fa926(p2281,p2285,p2287,p2314,p2315);
FA fa927(p2291,p2293,p2295,p2316,p2317);
HA ha231(p2297,p2299,p2318,p2319);
FA fa928(p2301,p2305,p2170,p2320,p2321);
FA fa929(p2172,p2176,p2178,p2322,p2323);
FA fa930(p2180,p2182,p2184,p2324,p2325);
FA fa931(p2190,p2196,p2198,p2326,p2327);
FA fa932(p2200,p2202,p2208,p2328,p2329);
HA ha232(p2212,p2307,p2330,p2331);
FA fa933(p2309,p2311,p2319,p2332,p2333);
FA fa934(p2204,p2206,p2224,p2334,p2335);
FA fa935(p2228,p2313,p2315,p2336,p2337);
FA fa936(p2317,p2321,p2331,p2338,p2339);
HA ha233(p2210,p2214,p2340,p2341);
FA fa937(p2216,p2232,p2323,p2342,p2343);
FA fa938(p2325,p2327,p2329,p2344,p2345);
FA fa939(p2333,p2218,p2220,p2346,p2347);
FA fa940(p2222,p2226,p2230,p2348,p2349);
FA fa941(p2236,p2335,p2337,p2350,p2351);
FA fa942(p2339,p2341,p2234,p2352,p2353);
FA fa943(p2343,p2345,p2238,p2354,p2355);
FA fa944(p2240,p2242,p2347,p2356,p2357);
FA fa945(p2349,p2351,p2353,p2358,p2359);
FA fa946(p2244,p2246,p2355,p2360,p2361);
HA ha234(p2248,p2250,p2362,p2363);
FA fa947(p2357,p2359,p2252,p2364,p2365);
FA fa948(p2254,p2361,p2363,p2366,p2367);
FA fa949(p2256,p2258,p2365,p2368,p2369);
FA fa950(p2260,p2367,p2262,p2370,p2371);
FA fa951(p2369,p2264,p2371,p2372,p2373);
FA fa952(p2266,p2373,p2268,p2374,p2375);
FA fa953(p2270,p2375,p2272,p2376,p2377);
HA ha235(ip_0_46,ip_1_45,p2378,p2379);
FA fa954(ip_2_44,ip_3_43,ip_4_42,p2380,p2381);
FA fa955(ip_5_41,ip_6_40,ip_7_39,p2382,p2383);
FA fa956(ip_8_38,ip_9_37,ip_10_36,p2384,p2385);
FA fa957(ip_11_35,ip_12_34,ip_13_33,p2386,p2387);
FA fa958(ip_14_32,ip_15_31,ip_16_30,p2388,p2389);
FA fa959(ip_17_29,ip_18_28,ip_19_27,p2390,p2391);
HA ha236(ip_20_26,ip_21_25,p2392,p2393);
FA fa960(ip_22_24,ip_23_23,ip_24_22,p2394,p2395);
FA fa961(ip_25_21,ip_26_20,ip_27_19,p2396,p2397);
FA fa962(ip_28_18,ip_29_17,ip_30_16,p2398,p2399);
FA fa963(ip_31_15,ip_32_14,ip_33_13,p2400,p2401);
HA ha237(ip_34_12,ip_35_11,p2402,p2403);
FA fa964(ip_36_10,ip_37_9,ip_38_8,p2404,p2405);
FA fa965(ip_39_7,ip_40_6,ip_41_5,p2406,p2407);
HA ha238(ip_42_4,ip_43_3,p2408,p2409);
FA fa966(ip_44_2,ip_45_1,ip_46_0,p2410,p2411);
FA fa967(p2282,p2288,p2302,p2412,p2413);
FA fa968(p2379,p2393,p2403,p2414,p2415);
HA ha239(p2409,p2381,p2416,p2417);
FA fa969(p2383,p2385,p2387,p2418,p2419);
FA fa970(p2389,p2391,p2395,p2420,p2421);
HA ha240(p2397,p2399,p2422,p2423);
HA ha241(p2401,p2405,p2424,p2425);
HA ha242(p2407,p2411,p2426,p2427);
FA fa971(p2274,p2276,p2278,p2428,p2429);
FA fa972(p2280,p2284,p2286,p2430,p2431);
FA fa973(p2290,p2292,p2294,p2432,p2433);
HA ha243(p2296,p2298,p2434,p2435);
HA ha244(p2300,p2304,p2436,p2437);
FA fa974(p2318,p2413,p2415,p2438,p2439);
FA fa975(p2417,p2423,p2425,p2440,p2441);
HA ha245(p2427,p2306,p2442,p2443);
FA fa976(p2308,p2310,p2330,p2444,p2445);
FA fa977(p2419,p2421,p2435,p2446,p2447);
FA fa978(p2437,p2312,p2314,p2448,p2449);
FA fa979(p2316,p2320,p2429,p2450,p2451);
FA fa980(p2431,p2433,p2439,p2452,p2453);
FA fa981(p2441,p2443,p2322,p2454,p2455);
FA fa982(p2324,p2326,p2328,p2456,p2457);
FA fa983(p2332,p2340,p2445,p2458,p2459);
HA ha246(p2447,p2334,p2460,p2461);
FA fa984(p2336,p2338,p2449,p2462,p2463);
FA fa985(p2451,p2453,p2455,p2464,p2465);
FA fa986(p2342,p2344,p2457,p2466,p2467);
FA fa987(p2459,p2461,p2346,p2468,p2469);
FA fa988(p2348,p2350,p2352,p2470,p2471);
HA ha247(p2463,p2465,p2472,p2473);
HA ha248(p2354,p2467,p2474,p2475);
FA fa989(p2469,p2473,p2356,p2476,p2477);
FA fa990(p2358,p2362,p2471,p2478,p2479);
FA fa991(p2475,p2360,p2477,p2480,p2481);
FA fa992(p2364,p2479,p2366,p2482,p2483);
HA ha249(p2481,p2368,p2484,p2485);
FA fa993(p2483,p2370,p2485,p2486,p2487);
FA fa994(p2372,p2487,p2374,p2488,p2489);
FA fa995(ip_0_47,ip_1_46,ip_2_45,p2490,p2491);
FA fa996(ip_3_44,ip_4_43,ip_5_42,p2492,p2493);
FA fa997(ip_6_41,ip_7_40,ip_8_39,p2494,p2495);
FA fa998(ip_9_38,ip_10_37,ip_11_36,p2496,p2497);
FA fa999(ip_12_35,ip_13_34,ip_14_33,p2498,p2499);
FA fa1000(ip_15_32,ip_16_31,ip_17_30,p2500,p2501);
FA fa1001(ip_18_29,ip_19_28,ip_20_27,p2502,p2503);
HA ha250(ip_21_26,ip_22_25,p2504,p2505);
FA fa1002(ip_23_24,ip_24_23,ip_25_22,p2506,p2507);
FA fa1003(ip_26_21,ip_27_20,ip_28_19,p2508,p2509);
FA fa1004(ip_29_18,ip_30_17,ip_31_16,p2510,p2511);
FA fa1005(ip_32_15,ip_33_14,ip_34_13,p2512,p2513);
FA fa1006(ip_35_12,ip_36_11,ip_37_10,p2514,p2515);
FA fa1007(ip_38_9,ip_39_8,ip_40_7,p2516,p2517);
FA fa1008(ip_41_6,ip_42_5,ip_43_4,p2518,p2519);
FA fa1009(ip_44_3,ip_45_2,ip_46_1,p2520,p2521);
HA ha251(ip_47_0,p2378,p2522,p2523);
HA ha252(p2392,p2402,p2524,p2525);
HA ha253(p2408,p2505,p2526,p2527);
FA fa1010(p2491,p2493,p2495,p2528,p2529);
FA fa1011(p2497,p2499,p2501,p2530,p2531);
FA fa1012(p2503,p2507,p2509,p2532,p2533);
FA fa1013(p2511,p2513,p2515,p2534,p2535);
FA fa1014(p2517,p2519,p2521,p2536,p2537);
FA fa1015(p2523,p2525,p2527,p2538,p2539);
FA fa1016(p2380,p2382,p2384,p2540,p2541);
FA fa1017(p2386,p2388,p2390,p2542,p2543);
FA fa1018(p2394,p2396,p2398,p2544,p2545);
FA fa1019(p2400,p2404,p2406,p2546,p2547);
FA fa1020(p2410,p2416,p2422,p2548,p2549);
FA fa1021(p2424,p2426,p2412,p2550,p2551);
FA fa1022(p2414,p2434,p2436,p2552,p2553);
FA fa1023(p2529,p2531,p2533,p2554,p2555);
HA ha254(p2535,p2537,p2556,p2557);
FA fa1024(p2539,p2418,p2420,p2558,p2559);
FA fa1025(p2442,p2541,p2543,p2560,p2561);
FA fa1026(p2545,p2547,p2549,p2562,p2563);
FA fa1027(p2551,p2557,p2428,p2564,p2565);
FA fa1028(p2430,p2432,p2438,p2566,p2567);
FA fa1029(p2440,p2553,p2555,p2568,p2569);
FA fa1030(p2444,p2446,p2559,p2570,p2571);
FA fa1031(p2561,p2563,p2565,p2572,p2573);
FA fa1032(p2448,p2450,p2452,p2574,p2575);
FA fa1033(p2454,p2460,p2567,p2576,p2577);
HA ha255(p2569,p2456,p2578,p2579);
FA fa1034(p2458,p2571,p2573,p2580,p2581);
FA fa1035(p2462,p2464,p2472,p2582,p2583);
FA fa1036(p2575,p2577,p2579,p2584,p2585);
FA fa1037(p2466,p2468,p2474,p2586,p2587);
FA fa1038(p2581,p2470,p2583,p2588,p2589);
FA fa1039(p2585,p2476,p2587,p2590,p2591);
FA fa1040(p2478,p2589,p2480,p2592,p2593);
FA fa1041(p2591,p2482,p2484,p2594,p2595);
FA fa1042(p2593,p2595,p2486,p2596,p2597);
FA fa1043(ip_0_48,ip_1_47,ip_2_46,p2598,p2599);
FA fa1044(ip_3_45,ip_4_44,ip_5_43,p2600,p2601);
HA ha256(ip_6_42,ip_7_41,p2602,p2603);
FA fa1045(ip_8_40,ip_9_39,ip_10_38,p2604,p2605);
HA ha257(ip_11_37,ip_12_36,p2606,p2607);
FA fa1046(ip_13_35,ip_14_34,ip_15_33,p2608,p2609);
FA fa1047(ip_16_32,ip_17_31,ip_18_30,p2610,p2611);
HA ha258(ip_19_29,ip_20_28,p2612,p2613);
FA fa1048(ip_21_27,ip_22_26,ip_23_25,p2614,p2615);
FA fa1049(ip_24_24,ip_25_23,ip_26_22,p2616,p2617);
FA fa1050(ip_27_21,ip_28_20,ip_29_19,p2618,p2619);
FA fa1051(ip_30_18,ip_31_17,ip_32_16,p2620,p2621);
FA fa1052(ip_33_15,ip_34_14,ip_35_13,p2622,p2623);
HA ha259(ip_36_12,ip_37_11,p2624,p2625);
FA fa1053(ip_38_10,ip_39_9,ip_40_8,p2626,p2627);
FA fa1054(ip_41_7,ip_42_6,ip_43_5,p2628,p2629);
FA fa1055(ip_44_4,ip_45_3,ip_46_2,p2630,p2631);
FA fa1056(ip_47_1,ip_48_0,p2504,p2632,p2633);
HA ha260(p2603,p2607,p2634,p2635);
HA ha261(p2613,p2625,p2636,p2637);
HA ha262(p2522,p2524,p2638,p2639);
HA ha263(p2526,p2599,p2640,p2641);
FA fa1057(p2601,p2605,p2609,p2642,p2643);
FA fa1058(p2611,p2615,p2617,p2644,p2645);
FA fa1059(p2619,p2621,p2623,p2646,p2647);
FA fa1060(p2627,p2629,p2631,p2648,p2649);
HA ha264(p2633,p2635,p2650,p2651);
FA fa1061(p2637,p2490,p2492,p2652,p2653);
FA fa1062(p2494,p2496,p2498,p2654,p2655);
FA fa1063(p2500,p2502,p2506,p2656,p2657);
FA fa1064(p2508,p2510,p2512,p2658,p2659);
FA fa1065(p2514,p2516,p2518,p2660,p2661);
FA fa1066(p2520,p2639,p2641,p2662,p2663);
FA fa1067(p2651,p2643,p2645,p2664,p2665);
FA fa1068(p2647,p2649,p2528,p2666,p2667);
FA fa1069(p2530,p2532,p2534,p2668,p2669);
FA fa1070(p2536,p2538,p2556,p2670,p2671);
FA fa1071(p2653,p2655,p2657,p2672,p2673);
HA ha265(p2659,p2661,p2674,p2675);
FA fa1072(p2663,p2540,p2542,p2676,p2677);
FA fa1073(p2544,p2546,p2548,p2678,p2679);
FA fa1074(p2550,p2665,p2667,p2680,p2681);
FA fa1075(p2675,p2552,p2554,p2682,p2683);
FA fa1076(p2669,p2671,p2673,p2684,p2685);
FA fa1077(p2558,p2560,p2562,p2686,p2687);
FA fa1078(p2564,p2677,p2679,p2688,p2689);
FA fa1079(p2681,p2566,p2568,p2690,p2691);
FA fa1080(p2683,p2685,p2570,p2692,p2693);
FA fa1081(p2572,p2578,p2687,p2694,p2695);
HA ha266(p2689,p2574,p2696,p2697);
FA fa1082(p2576,p2691,p2693,p2698,p2699);
FA fa1083(p2580,p2695,p2697,p2700,p2701);
FA fa1084(p2582,p2584,p2699,p2702,p2703);
FA fa1085(p2586,p2701,p2588,p2704,p2705);
HA ha267(p2703,p2590,p2706,p2707);
FA fa1086(p2705,p2592,p2707,p2708,p2709);
FA fa1087(p2594,p2709,p2596,p2710,p2711);
FA fa1088(ip_0_49,ip_1_48,ip_2_47,p2712,p2713);
FA fa1089(ip_3_46,ip_4_45,ip_5_44,p2714,p2715);
FA fa1090(ip_6_43,ip_7_42,ip_8_41,p2716,p2717);
FA fa1091(ip_9_40,ip_10_39,ip_11_38,p2718,p2719);
FA fa1092(ip_12_37,ip_13_36,ip_14_35,p2720,p2721);
FA fa1093(ip_15_34,ip_16_33,ip_17_32,p2722,p2723);
FA fa1094(ip_18_31,ip_19_30,ip_20_29,p2724,p2725);
FA fa1095(ip_21_28,ip_22_27,ip_23_26,p2726,p2727);
HA ha268(ip_24_25,ip_25_24,p2728,p2729);
FA fa1096(ip_26_23,ip_27_22,ip_28_21,p2730,p2731);
FA fa1097(ip_29_20,ip_30_19,ip_31_18,p2732,p2733);
HA ha269(ip_32_17,ip_33_16,p2734,p2735);
FA fa1098(ip_34_15,ip_35_14,ip_36_13,p2736,p2737);
HA ha270(ip_37_12,ip_38_11,p2738,p2739);
FA fa1099(ip_39_10,ip_40_9,ip_41_8,p2740,p2741);
HA ha271(ip_42_7,ip_43_6,p2742,p2743);
FA fa1100(ip_44_5,ip_45_4,ip_46_3,p2744,p2745);
HA ha272(ip_47_2,ip_48_1,p2746,p2747);
FA fa1101(ip_49_0,p2602,p2606,p2748,p2749);
FA fa1102(p2612,p2624,p2729,p2750,p2751);
FA fa1103(p2735,p2739,p2743,p2752,p2753);
FA fa1104(p2747,p2634,p2636,p2754,p2755);
FA fa1105(p2713,p2715,p2717,p2756,p2757);
FA fa1106(p2719,p2721,p2723,p2758,p2759);
FA fa1107(p2725,p2727,p2731,p2760,p2761);
FA fa1108(p2733,p2737,p2741,p2762,p2763);
FA fa1109(p2745,p2598,p2600,p2764,p2765);
HA ha273(p2604,p2608,p2766,p2767);
HA ha274(p2610,p2614,p2768,p2769);
FA fa1110(p2616,p2618,p2620,p2770,p2771);
FA fa1111(p2622,p2626,p2628,p2772,p2773);
FA fa1112(p2630,p2632,p2638,p2774,p2775);
HA ha275(p2640,p2650,p2776,p2777);
FA fa1113(p2749,p2751,p2753,p2778,p2779);
FA fa1114(p2755,p2757,p2759,p2780,p2781);
FA fa1115(p2761,p2763,p2767,p2782,p2783);
HA ha276(p2769,p2777,p2784,p2785);
FA fa1116(p2642,p2644,p2646,p2786,p2787);
FA fa1117(p2648,p2765,p2771,p2788,p2789);
FA fa1118(p2773,p2775,p2779,p2790,p2791);
FA fa1119(p2785,p2652,p2654,p2792,p2793);
FA fa1120(p2656,p2658,p2660,p2794,p2795);
FA fa1121(p2662,p2674,p2781,p2796,p2797);
FA fa1122(p2783,p2664,p2666,p2798,p2799);
FA fa1123(p2787,p2789,p2791,p2800,p2801);
FA fa1124(p2668,p2670,p2672,p2802,p2803);
FA fa1125(p2793,p2795,p2797,p2804,p2805);
FA fa1126(p2676,p2678,p2680,p2806,p2807);
FA fa1127(p2799,p2801,p2682,p2808,p2809);
FA fa1128(p2684,p2803,p2805,p2810,p2811);
HA ha277(p2686,p2688,p2812,p2813);
FA fa1129(p2807,p2809,p2690,p2814,p2815);
FA fa1130(p2692,p2696,p2811,p2816,p2817);
FA fa1131(p2813,p2694,p2815,p2818,p2819);
FA fa1132(p2698,p2817,p2700,p2820,p2821);
FA fa1133(p2819,p2702,p2821,p2822,p2823);
FA fa1134(p2704,p2706,p2823,p2824,p2825);
FA fa1135(p2825,p2708,p2710,p2826,p2827);
FA fa1136(ip_0_50,ip_1_49,ip_2_48,p2828,p2829);
FA fa1137(ip_3_47,ip_4_46,ip_5_45,p2830,p2831);
FA fa1138(ip_6_44,ip_7_43,ip_8_42,p2832,p2833);
HA ha278(ip_9_41,ip_10_40,p2834,p2835);
HA ha279(ip_11_39,ip_12_38,p2836,p2837);
FA fa1139(ip_13_37,ip_14_36,ip_15_35,p2838,p2839);
FA fa1140(ip_16_34,ip_17_33,ip_18_32,p2840,p2841);
FA fa1141(ip_19_31,ip_20_30,ip_21_29,p2842,p2843);
HA ha280(ip_22_28,ip_23_27,p2844,p2845);
FA fa1142(ip_24_26,ip_25_25,ip_26_24,p2846,p2847);
FA fa1143(ip_27_23,ip_28_22,ip_29_21,p2848,p2849);
FA fa1144(ip_30_20,ip_31_19,ip_32_18,p2850,p2851);
FA fa1145(ip_33_17,ip_34_16,ip_35_15,p2852,p2853);
FA fa1146(ip_36_14,ip_37_13,ip_38_12,p2854,p2855);
FA fa1147(ip_39_11,ip_40_10,ip_41_9,p2856,p2857);
FA fa1148(ip_42_8,ip_43_7,ip_44_6,p2858,p2859);
FA fa1149(ip_45_5,ip_46_4,ip_47_3,p2860,p2861);
FA fa1150(ip_48_2,ip_49_1,ip_50_0,p2862,p2863);
FA fa1151(p2728,p2734,p2738,p2864,p2865);
FA fa1152(p2742,p2746,p2835,p2866,p2867);
HA ha281(p2837,p2845,p2868,p2869);
FA fa1153(p2829,p2831,p2833,p2870,p2871);
FA fa1154(p2839,p2841,p2843,p2872,p2873);
FA fa1155(p2847,p2849,p2851,p2874,p2875);
FA fa1156(p2853,p2855,p2857,p2876,p2877);
FA fa1157(p2859,p2861,p2863,p2878,p2879);
FA fa1158(p2869,p2712,p2714,p2880,p2881);
FA fa1159(p2716,p2718,p2720,p2882,p2883);
HA ha282(p2722,p2724,p2884,p2885);
HA ha283(p2726,p2730,p2886,p2887);
HA ha284(p2732,p2736,p2888,p2889);
FA fa1160(p2740,p2744,p2865,p2890,p2891);
HA ha285(p2867,p2748,p2892,p2893);
FA fa1161(p2750,p2752,p2766,p2894,p2895);
FA fa1162(p2768,p2776,p2871,p2896,p2897);
FA fa1163(p2873,p2875,p2877,p2898,p2899);
HA ha286(p2879,p2885,p2900,p2901);
HA ha287(p2887,p2889,p2902,p2903);
FA fa1164(p2754,p2756,p2758,p2904,p2905);
FA fa1165(p2760,p2762,p2784,p2906,p2907);
FA fa1166(p2881,p2883,p2891,p2908,p2909);
HA ha288(p2893,p2901,p2910,p2911);
HA ha289(p2903,p2764,p2912,p2913);
FA fa1167(p2770,p2772,p2774,p2914,p2915);
FA fa1168(p2778,p2895,p2897,p2916,p2917);
FA fa1169(p2899,p2911,p2780,p2918,p2919);
FA fa1170(p2782,p2905,p2907,p2920,p2921);
FA fa1171(p2909,p2913,p2786,p2922,p2923);
FA fa1172(p2788,p2790,p2915,p2924,p2925);
HA ha290(p2917,p2919,p2926,p2927);
FA fa1173(p2792,p2794,p2796,p2928,p2929);
FA fa1174(p2921,p2923,p2927,p2930,p2931);
FA fa1175(p2798,p2800,p2925,p2932,p2933);
FA fa1176(p2802,p2804,p2929,p2934,p2935);
FA fa1177(p2931,p2806,p2808,p2936,p2937);
FA fa1178(p2812,p2933,p2810,p2938,p2939);
FA fa1179(p2935,p2814,p2937,p2940,p2941);
FA fa1180(p2939,p2816,p2818,p2942,p2943);
FA fa1181(p2941,p2820,p2943,p2944,p2945);
HA ha291(p2822,p2945,p2946,p2947);
FA fa1182(p2824,p2947,p2826,p2948,p2949);
FA fa1183(ip_0_51,ip_1_50,ip_2_49,p2950,p2951);
FA fa1184(ip_3_48,ip_4_47,ip_5_46,p2952,p2953);
FA fa1185(ip_6_45,ip_7_44,ip_8_43,p2954,p2955);
FA fa1186(ip_9_42,ip_10_41,ip_11_40,p2956,p2957);
FA fa1187(ip_12_39,ip_13_38,ip_14_37,p2958,p2959);
FA fa1188(ip_15_36,ip_16_35,ip_17_34,p2960,p2961);
FA fa1189(ip_18_33,ip_19_32,ip_20_31,p2962,p2963);
FA fa1190(ip_21_30,ip_22_29,ip_23_28,p2964,p2965);
FA fa1191(ip_24_27,ip_25_26,ip_26_25,p2966,p2967);
FA fa1192(ip_27_24,ip_28_23,ip_29_22,p2968,p2969);
FA fa1193(ip_30_21,ip_31_20,ip_32_19,p2970,p2971);
FA fa1194(ip_33_18,ip_34_17,ip_35_16,p2972,p2973);
FA fa1195(ip_36_15,ip_37_14,ip_38_13,p2974,p2975);
FA fa1196(ip_39_12,ip_40_11,ip_41_10,p2976,p2977);
FA fa1197(ip_42_9,ip_43_8,ip_44_7,p2978,p2979);
FA fa1198(ip_45_6,ip_46_5,ip_47_4,p2980,p2981);
FA fa1199(ip_48_3,ip_49_2,ip_50_1,p2982,p2983);
FA fa1200(ip_51_0,p2834,p2836,p2984,p2985);
FA fa1201(p2844,p2868,p2951,p2986,p2987);
FA fa1202(p2953,p2955,p2957,p2988,p2989);
FA fa1203(p2959,p2961,p2963,p2990,p2991);
FA fa1204(p2965,p2967,p2969,p2992,p2993);
FA fa1205(p2971,p2973,p2975,p2994,p2995);
FA fa1206(p2977,p2979,p2981,p2996,p2997);
FA fa1207(p2983,p2828,p2830,p2998,p2999);
FA fa1208(p2832,p2838,p2840,p3000,p3001);
FA fa1209(p2842,p2846,p2848,p3002,p3003);
FA fa1210(p2850,p2852,p2854,p3004,p3005);
FA fa1211(p2856,p2858,p2860,p3006,p3007);
FA fa1212(p2862,p2985,p2864,p3008,p3009);
FA fa1213(p2866,p2884,p2886,p3010,p3011);
HA ha292(p2888,p2987,p3012,p3013);
HA ha293(p2989,p2991,p3014,p3015);
FA fa1214(p2993,p2995,p2997,p3016,p3017);
FA fa1215(p2870,p2872,p2874,p3018,p3019);
FA fa1216(p2876,p2878,p2892,p3020,p3021);
FA fa1217(p2900,p2902,p2999,p3022,p3023);
FA fa1218(p3001,p3003,p3005,p3024,p3025);
FA fa1219(p3007,p3009,p3013,p3026,p3027);
FA fa1220(p3015,p2880,p2882,p3028,p3029);
FA fa1221(p2890,p2910,p3011,p3030,p3031);
FA fa1222(p3017,p2894,p2896,p3032,p3033);
FA fa1223(p2898,p2912,p3019,p3034,p3035);
FA fa1224(p3021,p3023,p3025,p3036,p3037);
FA fa1225(p3027,p2904,p2906,p3038,p3039);
FA fa1226(p2908,p3029,p3031,p3040,p3041);
HA ha294(p2914,p2916,p3042,p3043);
HA ha295(p2918,p2926,p3044,p3045);
FA fa1227(p3033,p3035,p3037,p3046,p3047);
FA fa1228(p2920,p2922,p3039,p3048,p3049);
FA fa1229(p3041,p3043,p3045,p3050,p3051);
FA fa1230(p2924,p3047,p2928,p3052,p3053);
FA fa1231(p2930,p3049,p3051,p3054,p3055);
FA fa1232(p2932,p3053,p2934,p3056,p3057);
FA fa1233(p3055,p2936,p2938,p3058,p3059);
FA fa1234(p3057,p2940,p3059,p3060,p3061);
FA fa1235(p2942,p3061,p2944,p3062,p3063);
FA fa1236(p2946,p3063,p2948,p3064,p3065);
FA fa1237(ip_0_52,ip_1_51,ip_2_50,p3066,p3067);
FA fa1238(ip_3_49,ip_4_48,ip_5_47,p3068,p3069);
FA fa1239(ip_6_46,ip_7_45,ip_8_44,p3070,p3071);
FA fa1240(ip_9_43,ip_10_42,ip_11_41,p3072,p3073);
FA fa1241(ip_12_40,ip_13_39,ip_14_38,p3074,p3075);
FA fa1242(ip_15_37,ip_16_36,ip_17_35,p3076,p3077);
FA fa1243(ip_18_34,ip_19_33,ip_20_32,p3078,p3079);
FA fa1244(ip_21_31,ip_22_30,ip_23_29,p3080,p3081);
HA ha296(ip_24_28,ip_25_27,p3082,p3083);
FA fa1245(ip_26_26,ip_27_25,ip_28_24,p3084,p3085);
FA fa1246(ip_29_23,ip_30_22,ip_31_21,p3086,p3087);
FA fa1247(ip_32_20,ip_33_19,ip_34_18,p3088,p3089);
HA ha297(ip_35_17,ip_36_16,p3090,p3091);
FA fa1248(ip_37_15,ip_38_14,ip_39_13,p3092,p3093);
FA fa1249(ip_40_12,ip_41_11,ip_42_10,p3094,p3095);
FA fa1250(ip_43_9,ip_44_8,ip_45_7,p3096,p3097);
FA fa1251(ip_46_6,ip_47_5,ip_48_4,p3098,p3099);
FA fa1252(ip_49_3,ip_50_2,ip_51_1,p3100,p3101);
FA fa1253(ip_52_0,p3083,p3091,p3102,p3103);
FA fa1254(p3067,p3069,p3071,p3104,p3105);
FA fa1255(p3073,p3075,p3077,p3106,p3107);
FA fa1256(p3079,p3081,p3085,p3108,p3109);
FA fa1257(p3087,p3089,p3093,p3110,p3111);
FA fa1258(p3095,p3097,p3099,p3112,p3113);
FA fa1259(p3101,p2950,p2952,p3114,p3115);
HA ha298(p2954,p2956,p3116,p3117);
FA fa1260(p2958,p2960,p2962,p3118,p3119);
FA fa1261(p2964,p2966,p2968,p3120,p3121);
FA fa1262(p2970,p2972,p2974,p3122,p3123);
FA fa1263(p2976,p2978,p2980,p3124,p3125);
FA fa1264(p2982,p3103,p2984,p3126,p3127);
FA fa1265(p3105,p3107,p3109,p3128,p3129);
FA fa1266(p3111,p3113,p3117,p3130,p3131);
FA fa1267(p2986,p2988,p2990,p3132,p3133);
FA fa1268(p2992,p2994,p2996,p3134,p3135);
FA fa1269(p3012,p3014,p3115,p3136,p3137);
FA fa1270(p3119,p3121,p3123,p3138,p3139);
FA fa1271(p3125,p3127,p2998,p3140,p3141);
FA fa1272(p3000,p3002,p3004,p3142,p3143);
FA fa1273(p3006,p3008,p3129,p3144,p3145);
FA fa1274(p3131,p3010,p3016,p3146,p3147);
FA fa1275(p3133,p3135,p3137,p3148,p3149);
HA ha299(p3139,p3141,p3150,p3151);
FA fa1276(p3018,p3020,p3022,p3152,p3153);
FA fa1277(p3024,p3026,p3143,p3154,p3155);
FA fa1278(p3145,p3151,p3028,p3156,p3157);
HA ha300(p3030,p3147,p3158,p3159);
FA fa1279(p3149,p3032,p3034,p3160,p3161);
FA fa1280(p3036,p3042,p3044,p3162,p3163);
FA fa1281(p3153,p3155,p3157,p3164,p3165);
FA fa1282(p3159,p3038,p3040,p3166,p3167);
HA ha301(p3046,p3161,p3168,p3169);
HA ha302(p3163,p3165,p3170,p3171);
FA fa1283(p3048,p3050,p3167,p3172,p3173);
FA fa1284(p3169,p3171,p3052,p3174,p3175);
HA ha303(p3054,p3173,p3176,p3177);
FA fa1285(p3175,p3056,p3177,p3178,p3179);
HA ha304(p3058,p3179,p3180,p3181);
FA fa1286(p3181,p3060,p3062,p3182,p3183);
FA fa1287(ip_0_53,ip_1_52,ip_2_51,p3184,p3185);
FA fa1288(ip_3_50,ip_4_49,ip_5_48,p3186,p3187);
HA ha305(ip_6_47,ip_7_46,p3188,p3189);
FA fa1289(ip_8_45,ip_9_44,ip_10_43,p3190,p3191);
FA fa1290(ip_11_42,ip_12_41,ip_13_40,p3192,p3193);
FA fa1291(ip_14_39,ip_15_38,ip_16_37,p3194,p3195);
FA fa1292(ip_17_36,ip_18_35,ip_19_34,p3196,p3197);
FA fa1293(ip_20_33,ip_21_32,ip_22_31,p3198,p3199);
FA fa1294(ip_23_30,ip_24_29,ip_25_28,p3200,p3201);
FA fa1295(ip_26_27,ip_27_26,ip_28_25,p3202,p3203);
FA fa1296(ip_29_24,ip_30_23,ip_31_22,p3204,p3205);
FA fa1297(ip_32_21,ip_33_20,ip_34_19,p3206,p3207);
FA fa1298(ip_35_18,ip_36_17,ip_37_16,p3208,p3209);
FA fa1299(ip_38_15,ip_39_14,ip_40_13,p3210,p3211);
FA fa1300(ip_41_12,ip_42_11,ip_43_10,p3212,p3213);
FA fa1301(ip_44_9,ip_45_8,ip_46_7,p3214,p3215);
FA fa1302(ip_47_6,ip_48_5,ip_49_4,p3216,p3217);
FA fa1303(ip_50_3,ip_51_2,ip_52_1,p3218,p3219);
FA fa1304(ip_53_0,p3082,p3090,p3220,p3221);
HA ha306(p3189,p3185,p3222,p3223);
FA fa1305(p3187,p3191,p3193,p3224,p3225);
FA fa1306(p3195,p3197,p3199,p3226,p3227);
HA ha307(p3201,p3203,p3228,p3229);
HA ha308(p3205,p3207,p3230,p3231);
FA fa1307(p3209,p3211,p3213,p3232,p3233);
FA fa1308(p3215,p3217,p3219,p3234,p3235);
FA fa1309(p3066,p3068,p3070,p3236,p3237);
HA ha309(p3072,p3074,p3238,p3239);
FA fa1310(p3076,p3078,p3080,p3240,p3241);
FA fa1311(p3084,p3086,p3088,p3242,p3243);
FA fa1312(p3092,p3094,p3096,p3244,p3245);
HA ha310(p3098,p3100,p3246,p3247);
FA fa1313(p3221,p3223,p3229,p3248,p3249);
FA fa1314(p3231,p3102,p3116,p3250,p3251);
FA fa1315(p3225,p3227,p3233,p3252,p3253);
HA ha311(p3235,p3239,p3254,p3255);
FA fa1316(p3247,p3104,p3106,p3256,p3257);
FA fa1317(p3108,p3110,p3112,p3258,p3259);
FA fa1318(p3237,p3241,p3243,p3260,p3261);
FA fa1319(p3245,p3249,p3255,p3262,p3263);
FA fa1320(p3114,p3118,p3120,p3264,p3265);
FA fa1321(p3122,p3124,p3126,p3266,p3267);
FA fa1322(p3251,p3253,p3128,p3268,p3269);
FA fa1323(p3130,p3257,p3259,p3270,p3271);
FA fa1324(p3261,p3263,p3132,p3272,p3273);
FA fa1325(p3134,p3136,p3138,p3274,p3275);
HA ha312(p3140,p3150,p3276,p3277);
FA fa1326(p3265,p3267,p3269,p3278,p3279);
FA fa1327(p3142,p3144,p3271,p3280,p3281);
FA fa1328(p3273,p3277,p3146,p3282,p3283);
FA fa1329(p3148,p3158,p3275,p3284,p3285);
FA fa1330(p3279,p3152,p3154,p3286,p3287);
FA fa1331(p3156,p3281,p3283,p3288,p3289);
FA fa1332(p3285,p3160,p3162,p3290,p3291);
FA fa1333(p3164,p3168,p3170,p3292,p3293);
FA fa1334(p3287,p3289,p3166,p3294,p3295);
FA fa1335(p3291,p3293,p3295,p3296,p3297);
FA fa1336(p3172,p3174,p3176,p3298,p3299);
FA fa1337(p3297,p3299,p3178,p3300,p3301);
HA ha313(p3180,p3301,p3302,p3303);
FA fa1338(ip_0_54,ip_1_53,ip_2_52,p3304,p3305);
FA fa1339(ip_3_51,ip_4_50,ip_5_49,p3306,p3307);
FA fa1340(ip_6_48,ip_7_47,ip_8_46,p3308,p3309);
FA fa1341(ip_9_45,ip_10_44,ip_11_43,p3310,p3311);
FA fa1342(ip_12_42,ip_13_41,ip_14_40,p3312,p3313);
FA fa1343(ip_15_39,ip_16_38,ip_17_37,p3314,p3315);
HA ha314(ip_18_36,ip_19_35,p3316,p3317);
FA fa1344(ip_20_34,ip_21_33,ip_22_32,p3318,p3319);
FA fa1345(ip_23_31,ip_24_30,ip_25_29,p3320,p3321);
HA ha315(ip_26_28,ip_27_27,p3322,p3323);
FA fa1346(ip_28_26,ip_29_25,ip_30_24,p3324,p3325);
FA fa1347(ip_31_23,ip_32_22,ip_33_21,p3326,p3327);
FA fa1348(ip_34_20,ip_35_19,ip_36_18,p3328,p3329);
HA ha316(ip_37_17,ip_38_16,p3330,p3331);
FA fa1349(ip_39_15,ip_40_14,ip_41_13,p3332,p3333);
HA ha317(ip_42_12,ip_43_11,p3334,p3335);
FA fa1350(ip_44_10,ip_45_9,ip_46_8,p3336,p3337);
FA fa1351(ip_47_7,ip_48_6,ip_49_5,p3338,p3339);
FA fa1352(ip_50_4,ip_51_3,ip_52_2,p3340,p3341);
FA fa1353(ip_53_1,ip_54_0,p3188,p3342,p3343);
FA fa1354(p3317,p3323,p3331,p3344,p3345);
FA fa1355(p3335,p3305,p3307,p3346,p3347);
HA ha318(p3309,p3311,p3348,p3349);
HA ha319(p3313,p3315,p3350,p3351);
FA fa1356(p3319,p3321,p3325,p3352,p3353);
FA fa1357(p3327,p3329,p3333,p3354,p3355);
FA fa1358(p3337,p3339,p3341,p3356,p3357);
FA fa1359(p3343,p3184,p3186,p3358,p3359);
FA fa1360(p3190,p3192,p3194,p3360,p3361);
FA fa1361(p3196,p3198,p3200,p3362,p3363);
HA ha320(p3202,p3204,p3364,p3365);
FA fa1362(p3206,p3208,p3210,p3366,p3367);
FA fa1363(p3212,p3214,p3216,p3368,p3369);
FA fa1364(p3218,p3222,p3228,p3370,p3371);
FA fa1365(p3230,p3345,p3349,p3372,p3373);
FA fa1366(p3351,p3220,p3238,p3374,p3375);
FA fa1367(p3246,p3347,p3353,p3376,p3377);
HA ha321(p3355,p3357,p3378,p3379);
HA ha322(p3365,p3224,p3380,p3381);
FA fa1368(p3226,p3232,p3234,p3382,p3383);
FA fa1369(p3254,p3359,p3361,p3384,p3385);
FA fa1370(p3363,p3367,p3369,p3386,p3387);
FA fa1371(p3371,p3373,p3379,p3388,p3389);
FA fa1372(p3236,p3240,p3242,p3390,p3391);
HA ha323(p3244,p3248,p3392,p3393);
FA fa1373(p3375,p3377,p3381,p3394,p3395);
FA fa1374(p3250,p3252,p3383,p3396,p3397);
FA fa1375(p3385,p3387,p3389,p3398,p3399);
FA fa1376(p3393,p3256,p3258,p3400,p3401);
HA ha324(p3260,p3262,p3402,p3403);
HA ha325(p3391,p3395,p3404,p3405);
FA fa1377(p3264,p3266,p3268,p3406,p3407);
FA fa1378(p3276,p3397,p3399,p3408,p3409);
FA fa1379(p3403,p3405,p3270,p3410,p3411);
FA fa1380(p3272,p3401,p3274,p3412,p3413);
FA fa1381(p3278,p3407,p3409,p3414,p3415);
FA fa1382(p3411,p3280,p3282,p3416,p3417);
FA fa1383(p3413,p3284,p3415,p3418,p3419);
FA fa1384(p3286,p3288,p3417,p3420,p3421);
FA fa1385(p3419,p3290,p3292,p3422,p3423);
HA ha326(p3294,p3421,p3424,p3425);
FA fa1386(p3425,p3296,p3423,p3426,p3427);
FA fa1387(p3298,p3427,p3300,p3428,p3429);
FA fa1388(ip_0_55,ip_1_54,ip_2_53,p3430,p3431);
HA ha327(ip_3_52,ip_4_51,p3432,p3433);
FA fa1389(ip_5_50,ip_6_49,ip_7_48,p3434,p3435);
FA fa1390(ip_8_47,ip_9_46,ip_10_45,p3436,p3437);
FA fa1391(ip_11_44,ip_12_43,ip_13_42,p3438,p3439);
FA fa1392(ip_14_41,ip_15_40,ip_16_39,p3440,p3441);
FA fa1393(ip_17_38,ip_18_37,ip_19_36,p3442,p3443);
FA fa1394(ip_20_35,ip_21_34,ip_22_33,p3444,p3445);
FA fa1395(ip_23_32,ip_24_31,ip_25_30,p3446,p3447);
FA fa1396(ip_26_29,ip_27_28,ip_28_27,p3448,p3449);
FA fa1397(ip_29_26,ip_30_25,ip_31_24,p3450,p3451);
FA fa1398(ip_32_23,ip_33_22,ip_34_21,p3452,p3453);
FA fa1399(ip_35_20,ip_36_19,ip_37_18,p3454,p3455);
HA ha328(ip_38_17,ip_39_16,p3456,p3457);
FA fa1400(ip_40_15,ip_41_14,ip_42_13,p3458,p3459);
FA fa1401(ip_43_12,ip_44_11,ip_45_10,p3460,p3461);
FA fa1402(ip_46_9,ip_47_8,ip_48_7,p3462,p3463);
HA ha329(ip_49_6,ip_50_5,p3464,p3465);
FA fa1403(ip_51_4,ip_52_3,ip_53_2,p3466,p3467);
FA fa1404(ip_54_1,ip_55_0,p3316,p3468,p3469);
FA fa1405(p3322,p3330,p3334,p3470,p3471);
HA ha330(p3433,p3457,p3472,p3473);
FA fa1406(p3465,p3431,p3435,p3474,p3475);
HA ha331(p3437,p3439,p3476,p3477);
FA fa1407(p3441,p3443,p3445,p3478,p3479);
FA fa1408(p3447,p3449,p3451,p3480,p3481);
HA ha332(p3453,p3455,p3482,p3483);
FA fa1409(p3459,p3461,p3463,p3484,p3485);
FA fa1410(p3467,p3469,p3473,p3486,p3487);
FA fa1411(p3304,p3306,p3308,p3488,p3489);
FA fa1412(p3310,p3312,p3314,p3490,p3491);
HA ha333(p3318,p3320,p3492,p3493);
FA fa1413(p3324,p3326,p3328,p3494,p3495);
HA ha334(p3332,p3336,p3496,p3497);
FA fa1414(p3338,p3340,p3342,p3498,p3499);
FA fa1415(p3348,p3350,p3471,p3500,p3501);
FA fa1416(p3477,p3483,p3344,p3502,p3503);
FA fa1417(p3364,p3475,p3479,p3504,p3505);
FA fa1418(p3481,p3485,p3487,p3506,p3507);
FA fa1419(p3493,p3497,p3346,p3508,p3509);
FA fa1420(p3352,p3354,p3356,p3510,p3511);
FA fa1421(p3378,p3489,p3491,p3512,p3513);
FA fa1422(p3495,p3499,p3501,p3514,p3515);
HA ha335(p3503,p3358,p3516,p3517);
HA ha336(p3360,p3362,p3518,p3519);
FA fa1423(p3366,p3368,p3370,p3520,p3521);
FA fa1424(p3372,p3380,p3505,p3522,p3523);
FA fa1425(p3507,p3509,p3374,p3524,p3525);
HA ha337(p3376,p3392,p3526,p3527);
FA fa1426(p3511,p3513,p3515,p3528,p3529);
FA fa1427(p3517,p3519,p3382,p3530,p3531);
FA fa1428(p3384,p3386,p3388,p3532,p3533);
FA fa1429(p3521,p3523,p3525,p3534,p3535);
HA ha338(p3527,p3390,p3536,p3537);
HA ha339(p3394,p3402,p3538,p3539);
FA fa1430(p3404,p3529,p3531,p3540,p3541);
FA fa1431(p3396,p3398,p3533,p3542,p3543);
FA fa1432(p3535,p3537,p3539,p3544,p3545);
HA ha340(p3400,p3541,p3546,p3547);
FA fa1433(p3406,p3408,p3410,p3548,p3549);
FA fa1434(p3543,p3545,p3547,p3550,p3551);
FA fa1435(p3412,p3414,p3549,p3552,p3553);
FA fa1436(p3551,p3416,p3418,p3554,p3555);
FA fa1437(p3553,p3420,p3424,p3556,p3557);
FA fa1438(p3555,p3422,p3557,p3558,p3559);
FA fa1439(p3426,p3559,p3428,p3560,p3561);
FA fa1440(ip_0_56,ip_1_55,ip_2_54,p3562,p3563);
FA fa1441(ip_3_53,ip_4_52,ip_5_51,p3564,p3565);
FA fa1442(ip_6_50,ip_7_49,ip_8_48,p3566,p3567);
FA fa1443(ip_9_47,ip_10_46,ip_11_45,p3568,p3569);
HA ha341(ip_12_44,ip_13_43,p3570,p3571);
FA fa1444(ip_14_42,ip_15_41,ip_16_40,p3572,p3573);
FA fa1445(ip_17_39,ip_18_38,ip_19_37,p3574,p3575);
FA fa1446(ip_20_36,ip_21_35,ip_22_34,p3576,p3577);
FA fa1447(ip_23_33,ip_24_32,ip_25_31,p3578,p3579);
FA fa1448(ip_26_30,ip_27_29,ip_28_28,p3580,p3581);
FA fa1449(ip_29_27,ip_30_26,ip_31_25,p3582,p3583);
FA fa1450(ip_32_24,ip_33_23,ip_34_22,p3584,p3585);
FA fa1451(ip_35_21,ip_36_20,ip_37_19,p3586,p3587);
FA fa1452(ip_38_18,ip_39_17,ip_40_16,p3588,p3589);
FA fa1453(ip_41_15,ip_42_14,ip_43_13,p3590,p3591);
FA fa1454(ip_44_12,ip_45_11,ip_46_10,p3592,p3593);
HA ha342(ip_47_9,ip_48_8,p3594,p3595);
HA ha343(ip_49_7,ip_50_6,p3596,p3597);
FA fa1455(ip_51_5,ip_52_4,ip_53_3,p3598,p3599);
HA ha344(ip_54_2,ip_55_1,p3600,p3601);
FA fa1456(ip_56_0,p3432,p3456,p3602,p3603);
FA fa1457(p3464,p3571,p3595,p3604,p3605);
HA ha345(p3597,p3601,p3606,p3607);
FA fa1458(p3472,p3563,p3565,p3608,p3609);
FA fa1459(p3567,p3569,p3573,p3610,p3611);
FA fa1460(p3575,p3577,p3579,p3612,p3613);
FA fa1461(p3581,p3583,p3585,p3614,p3615);
FA fa1462(p3587,p3589,p3591,p3616,p3617);
FA fa1463(p3593,p3599,p3607,p3618,p3619);
FA fa1464(p3430,p3434,p3436,p3620,p3621);
HA ha346(p3438,p3440,p3622,p3623);
FA fa1465(p3442,p3444,p3446,p3624,p3625);
HA ha347(p3448,p3450,p3626,p3627);
FA fa1466(p3452,p3454,p3458,p3628,p3629);
FA fa1467(p3460,p3462,p3466,p3630,p3631);
FA fa1468(p3468,p3476,p3482,p3632,p3633);
HA ha348(p3603,p3605,p3634,p3635);
FA fa1469(p3470,p3492,p3496,p3636,p3637);
FA fa1470(p3609,p3611,p3613,p3638,p3639);
FA fa1471(p3615,p3617,p3619,p3640,p3641);
HA ha349(p3623,p3627,p3642,p3643);
FA fa1472(p3635,p3474,p3478,p3644,p3645);
HA ha350(p3480,p3484,p3646,p3647);
FA fa1473(p3486,p3621,p3625,p3648,p3649);
FA fa1474(p3629,p3631,p3633,p3650,p3651);
FA fa1475(p3643,p3488,p3490,p3652,p3653);
HA ha351(p3494,p3498,p3654,p3655);
FA fa1476(p3500,p3502,p3637,p3656,p3657);
FA fa1477(p3639,p3641,p3647,p3658,p3659);
FA fa1478(p3504,p3506,p3508,p3660,p3661);
FA fa1479(p3516,p3518,p3645,p3662,p3663);
FA fa1480(p3649,p3651,p3655,p3664,p3665);
HA ha352(p3510,p3512,p3666,p3667);
FA fa1481(p3514,p3526,p3653,p3668,p3669);
FA fa1482(p3657,p3659,p3520,p3670,p3671);
FA fa1483(p3522,p3524,p3661,p3672,p3673);
FA fa1484(p3663,p3665,p3667,p3674,p3675);
FA fa1485(p3528,p3530,p3536,p3676,p3677);
FA fa1486(p3538,p3669,p3671,p3678,p3679);
FA fa1487(p3532,p3534,p3673,p3680,p3681);
FA fa1488(p3675,p3540,p3546,p3682,p3683);
HA ha353(p3677,p3679,p3684,p3685);
HA ha354(p3542,p3544,p3686,p3687);
FA fa1489(p3681,p3685,p3683,p3688,p3689);
FA fa1490(p3687,p3548,p3550,p3690,p3691);
HA ha355(p3689,p3552,p3692,p3693);
HA ha356(p3691,p3554,p3694,p3695);
FA fa1491(p3693,p3695,p3556,p3696,p3697);
FA fa1492(p3697,p3558,p3560,p3698,p3699);
HA ha357(ip_0_57,ip_1_56,p3700,p3701);
FA fa1493(ip_2_55,ip_3_54,ip_4_53,p3702,p3703);
FA fa1494(ip_5_52,ip_6_51,ip_7_50,p3704,p3705);
HA ha358(ip_8_49,ip_9_48,p3706,p3707);
FA fa1495(ip_10_47,ip_11_46,ip_12_45,p3708,p3709);
FA fa1496(ip_13_44,ip_14_43,ip_15_42,p3710,p3711);
FA fa1497(ip_16_41,ip_17_40,ip_18_39,p3712,p3713);
FA fa1498(ip_19_38,ip_20_37,ip_21_36,p3714,p3715);
FA fa1499(ip_22_35,ip_23_34,ip_24_33,p3716,p3717);
FA fa1500(ip_25_32,ip_26_31,ip_27_30,p3718,p3719);
HA ha359(ip_28_29,ip_29_28,p3720,p3721);
FA fa1501(ip_30_27,ip_31_26,ip_32_25,p3722,p3723);
FA fa1502(ip_33_24,ip_34_23,ip_35_22,p3724,p3725);
FA fa1503(ip_36_21,ip_37_20,ip_38_19,p3726,p3727);
FA fa1504(ip_39_18,ip_40_17,ip_41_16,p3728,p3729);
FA fa1505(ip_42_15,ip_43_14,ip_44_13,p3730,p3731);
FA fa1506(ip_45_12,ip_46_11,ip_47_10,p3732,p3733);
FA fa1507(ip_48_9,ip_49_8,ip_50_7,p3734,p3735);
FA fa1508(ip_51_6,ip_52_5,ip_53_4,p3736,p3737);
FA fa1509(ip_54_3,ip_55_2,ip_56_1,p3738,p3739);
FA fa1510(ip_57_0,p3570,p3594,p3740,p3741);
FA fa1511(p3596,p3600,p3701,p3742,p3743);
FA fa1512(p3707,p3721,p3606,p3744,p3745);
FA fa1513(p3703,p3705,p3709,p3746,p3747);
FA fa1514(p3711,p3713,p3715,p3748,p3749);
HA ha360(p3717,p3719,p3750,p3751);
FA fa1515(p3723,p3725,p3727,p3752,p3753);
HA ha361(p3729,p3731,p3754,p3755);
FA fa1516(p3733,p3735,p3737,p3756,p3757);
FA fa1517(p3739,p3562,p3564,p3758,p3759);
HA ha362(p3566,p3568,p3760,p3761);
FA fa1518(p3572,p3574,p3576,p3762,p3763);
FA fa1519(p3578,p3580,p3582,p3764,p3765);
FA fa1520(p3584,p3586,p3588,p3766,p3767);
FA fa1521(p3590,p3592,p3598,p3768,p3769);
HA ha363(p3741,p3743,p3770,p3771);
FA fa1522(p3745,p3751,p3755,p3772,p3773);
FA fa1523(p3602,p3604,p3622,p3774,p3775);
FA fa1524(p3626,p3634,p3747,p3776,p3777);
FA fa1525(p3749,p3753,p3757,p3778,p3779);
HA ha364(p3761,p3771,p3780,p3781);
HA ha365(p3608,p3610,p3782,p3783);
FA fa1526(p3612,p3614,p3616,p3784,p3785);
FA fa1527(p3618,p3642,p3759,p3786,p3787);
FA fa1528(p3763,p3765,p3767,p3788,p3789);
FA fa1529(p3769,p3773,p3781,p3790,p3791);
FA fa1530(p3620,p3624,p3628,p3792,p3793);
FA fa1531(p3630,p3632,p3646,p3794,p3795);
FA fa1532(p3775,p3777,p3779,p3796,p3797);
HA ha366(p3783,p3636,p3798,p3799);
FA fa1533(p3638,p3640,p3654,p3800,p3801);
FA fa1534(p3785,p3787,p3789,p3802,p3803);
FA fa1535(p3791,p3644,p3648,p3804,p3805);
HA ha367(p3650,p3793,p3806,p3807);
FA fa1536(p3795,p3797,p3799,p3808,p3809);
FA fa1537(p3652,p3656,p3658,p3810,p3811);
HA ha368(p3666,p3801,p3812,p3813);
FA fa1538(p3803,p3807,p3660,p3814,p3815);
FA fa1539(p3662,p3664,p3805,p3816,p3817);
FA fa1540(p3809,p3813,p3668,p3818,p3819);
FA fa1541(p3670,p3811,p3815,p3820,p3821);
FA fa1542(p3672,p3674,p3817,p3822,p3823);
FA fa1543(p3819,p3676,p3678,p3824,p3825);
FA fa1544(p3684,p3821,p3680,p3826,p3827);
FA fa1545(p3686,p3823,p3682,p3828,p3829);
FA fa1546(p3825,p3827,p3688,p3830,p3831);
HA ha369(p3829,p3831,p3832,p3833);
FA fa1547(p3690,p3692,p3833,p3834,p3835);
HA ha370(p3694,p3835,p3836,p3837);
FA fa1548(p3837,p3696,p3698,p3838,p3839);
FA fa1549(ip_0_58,ip_1_57,ip_2_56,p3840,p3841);
FA fa1550(ip_3_55,ip_4_54,ip_5_53,p3842,p3843);
FA fa1551(ip_6_52,ip_7_51,ip_8_50,p3844,p3845);
HA ha371(ip_9_49,ip_10_48,p3846,p3847);
FA fa1552(ip_11_47,ip_12_46,ip_13_45,p3848,p3849);
HA ha372(ip_14_44,ip_15_43,p3850,p3851);
FA fa1553(ip_16_42,ip_17_41,ip_18_40,p3852,p3853);
FA fa1554(ip_19_39,ip_20_38,ip_21_37,p3854,p3855);
FA fa1555(ip_22_36,ip_23_35,ip_24_34,p3856,p3857);
FA fa1556(ip_25_33,ip_26_32,ip_27_31,p3858,p3859);
FA fa1557(ip_28_30,ip_29_29,ip_30_28,p3860,p3861);
HA ha373(ip_31_27,ip_32_26,p3862,p3863);
FA fa1558(ip_33_25,ip_34_24,ip_35_23,p3864,p3865);
FA fa1559(ip_36_22,ip_37_21,ip_38_20,p3866,p3867);
FA fa1560(ip_39_19,ip_40_18,ip_41_17,p3868,p3869);
FA fa1561(ip_42_16,ip_43_15,ip_44_14,p3870,p3871);
FA fa1562(ip_45_13,ip_46_12,ip_47_11,p3872,p3873);
HA ha374(ip_48_10,ip_49_9,p3874,p3875);
HA ha375(ip_50_8,ip_51_7,p3876,p3877);
FA fa1563(ip_52_6,ip_53_5,ip_54_4,p3878,p3879);
FA fa1564(ip_55_3,ip_56_2,ip_57_1,p3880,p3881);
FA fa1565(ip_58_0,p3700,p3706,p3882,p3883);
HA ha376(p3720,p3847,p3884,p3885);
FA fa1566(p3851,p3863,p3875,p3886,p3887);
FA fa1567(p3877,p3841,p3843,p3888,p3889);
HA ha377(p3845,p3849,p3890,p3891);
FA fa1568(p3853,p3855,p3857,p3892,p3893);
HA ha378(p3859,p3861,p3894,p3895);
FA fa1569(p3865,p3867,p3869,p3896,p3897);
FA fa1570(p3871,p3873,p3879,p3898,p3899);
FA fa1571(p3881,p3885,p3702,p3900,p3901);
HA ha379(p3704,p3708,p3902,p3903);
FA fa1572(p3710,p3712,p3714,p3904,p3905);
HA ha380(p3716,p3718,p3906,p3907);
HA ha381(p3722,p3724,p3908,p3909);
FA fa1573(p3726,p3728,p3730,p3910,p3911);
FA fa1574(p3732,p3734,p3736,p3912,p3913);
FA fa1575(p3738,p3750,p3754,p3914,p3915);
FA fa1576(p3883,p3887,p3891,p3916,p3917);
FA fa1577(p3895,p3740,p3742,p3918,p3919);
HA ha382(p3744,p3760,p3920,p3921);
FA fa1578(p3770,p3889,p3893,p3922,p3923);
FA fa1579(p3897,p3899,p3901,p3924,p3925);
FA fa1580(p3903,p3907,p3909,p3926,p3927);
FA fa1581(p3746,p3748,p3752,p3928,p3929);
FA fa1582(p3756,p3780,p3905,p3930,p3931);
FA fa1583(p3911,p3913,p3915,p3932,p3933);
HA ha383(p3917,p3921,p3934,p3935);
HA ha384(p3758,p3762,p3936,p3937);
FA fa1584(p3764,p3766,p3768,p3938,p3939);
FA fa1585(p3772,p3782,p3919,p3940,p3941);
HA ha385(p3923,p3925,p3942,p3943);
FA fa1586(p3927,p3935,p3774,p3944,p3945);
HA ha386(p3776,p3778,p3946,p3947);
FA fa1587(p3929,p3931,p3933,p3948,p3949);
FA fa1588(p3937,p3943,p3784,p3950,p3951);
FA fa1589(p3786,p3788,p3790,p3952,p3953);
FA fa1590(p3798,p3939,p3941,p3954,p3955);
FA fa1591(p3945,p3947,p3792,p3956,p3957);
FA fa1592(p3794,p3796,p3806,p3958,p3959);
HA ha387(p3949,p3951,p3960,p3961);
HA ha388(p3800,p3802,p3962,p3963);
FA fa1593(p3812,p3953,p3955,p3964,p3965);
FA fa1594(p3957,p3961,p3804,p3966,p3967);
FA fa1595(p3808,p3959,p3963,p3968,p3969);
HA ha389(p3810,p3814,p3970,p3971);
FA fa1596(p3965,p3967,p3816,p3972,p3973);
FA fa1597(p3818,p3969,p3971,p3974,p3975);
FA fa1598(p3820,p3973,p3822,p3976,p3977);
FA fa1599(p3975,p3824,p3826,p3978,p3979);
FA fa1600(p3977,p3828,p3830,p3980,p3981);
FA fa1601(p3832,p3979,p3981,p3982,p3983);
FA fa1602(p3983,p3834,p3836,p3984,p3985);
FA fa1603(ip_0_59,ip_1_58,ip_2_57,p3986,p3987);
FA fa1604(ip_3_56,ip_4_55,ip_5_54,p3988,p3989);
HA ha390(ip_6_53,ip_7_52,p3990,p3991);
FA fa1605(ip_8_51,ip_9_50,ip_10_49,p3992,p3993);
FA fa1606(ip_11_48,ip_12_47,ip_13_46,p3994,p3995);
FA fa1607(ip_14_45,ip_15_44,ip_16_43,p3996,p3997);
HA ha391(ip_17_42,ip_18_41,p3998,p3999);
FA fa1608(ip_19_40,ip_20_39,ip_21_38,p4000,p4001);
FA fa1609(ip_22_37,ip_23_36,ip_24_35,p4002,p4003);
FA fa1610(ip_25_34,ip_26_33,ip_27_32,p4004,p4005);
FA fa1611(ip_28_31,ip_29_30,ip_30_29,p4006,p4007);
FA fa1612(ip_31_28,ip_32_27,ip_33_26,p4008,p4009);
FA fa1613(ip_34_25,ip_35_24,ip_36_23,p4010,p4011);
HA ha392(ip_37_22,ip_38_21,p4012,p4013);
FA fa1614(ip_39_20,ip_40_19,ip_41_18,p4014,p4015);
FA fa1615(ip_42_17,ip_43_16,ip_44_15,p4016,p4017);
FA fa1616(ip_45_14,ip_46_13,ip_47_12,p4018,p4019);
FA fa1617(ip_48_11,ip_49_10,ip_50_9,p4020,p4021);
HA ha393(ip_51_8,ip_52_7,p4022,p4023);
HA ha394(ip_53_6,ip_54_5,p4024,p4025);
FA fa1618(ip_55_4,ip_56_3,ip_57_2,p4026,p4027);
FA fa1619(ip_58_1,ip_59_0,p3846,p4028,p4029);
HA ha395(p3850,p3862,p4030,p4031);
FA fa1620(p3874,p3876,p3991,p4032,p4033);
HA ha396(p3999,p4013,p4034,p4035);
FA fa1621(p4023,p4025,p3884,p4036,p4037);
FA fa1622(p3987,p3989,p3993,p4038,p4039);
FA fa1623(p3995,p3997,p4001,p4040,p4041);
FA fa1624(p4003,p4005,p4007,p4042,p4043);
FA fa1625(p4009,p4011,p4015,p4044,p4045);
FA fa1626(p4017,p4019,p4021,p4046,p4047);
FA fa1627(p4027,p4029,p4031,p4048,p4049);
FA fa1628(p4035,p3840,p3842,p4050,p4051);
HA ha397(p3844,p3848,p4052,p4053);
FA fa1629(p3852,p3854,p3856,p4054,p4055);
HA ha398(p3858,p3860,p4056,p4057);
FA fa1630(p3864,p3866,p3868,p4058,p4059);
FA fa1631(p3870,p3872,p3878,p4060,p4061);
FA fa1632(p3880,p3890,p3894,p4062,p4063);
FA fa1633(p4033,p4037,p3882,p4064,p4065);
HA ha399(p3886,p3902,p4066,p4067);
HA ha400(p3906,p3908,p4068,p4069);
HA ha401(p4039,p4041,p4070,p4071);
FA fa1634(p4043,p4045,p4047,p4072,p4073);
HA ha402(p4049,p4053,p4074,p4075);
FA fa1635(p4057,p3888,p3892,p4076,p4077);
HA ha403(p3896,p3898,p4078,p4079);
HA ha404(p3900,p3920,p4080,p4081);
HA ha405(p4051,p4055,p4082,p4083);
FA fa1636(p4059,p4061,p4063,p4084,p4085);
FA fa1637(p4065,p4067,p4069,p4086,p4087);
FA fa1638(p4071,p4075,p3904,p4088,p4089);
FA fa1639(p3910,p3912,p3914,p4090,p4091);
FA fa1640(p3916,p3934,p4073,p4092,p4093);
HA ha406(p4079,p4081,p4094,p4095);
FA fa1641(p4083,p3918,p3922,p4096,p4097);
FA fa1642(p3924,p3926,p3936,p4098,p4099);
FA fa1643(p3942,p4077,p4085,p4100,p4101);
FA fa1644(p4087,p4089,p4095,p4102,p4103);
FA fa1645(p3928,p3930,p3932,p4104,p4105);
FA fa1646(p3946,p4091,p4093,p4106,p4107);
FA fa1647(p3938,p3940,p3944,p4108,p4109);
FA fa1648(p4097,p4099,p4101,p4110,p4111);
FA fa1649(p4103,p3948,p3950,p4112,p4113);
FA fa1650(p3960,p4105,p4107,p4114,p4115);
FA fa1651(p3952,p3954,p3956,p4116,p4117);
FA fa1652(p3962,p4109,p4111,p4118,p4119);
FA fa1653(p3958,p4113,p4115,p4120,p4121);
FA fa1654(p3964,p3966,p3970,p4122,p4123);
FA fa1655(p4117,p4119,p3968,p4124,p4125);
FA fa1656(p4121,p3972,p4123,p4126,p4127);
FA fa1657(p4125,p3974,p3976,p4128,p4129);
FA fa1658(p4127,p4129,p3978,p4130,p4131);
HA ha407(p3980,p4131,p4132,p4133);
FA fa1659(p3982,p4133,p3984,p4134,p4135);
FA fa1660(ip_0_60,ip_1_59,ip_2_58,p4136,p4137);
FA fa1661(ip_3_57,ip_4_56,ip_5_55,p4138,p4139);
HA ha408(ip_6_54,ip_7_53,p4140,p4141);
FA fa1662(ip_8_52,ip_9_51,ip_10_50,p4142,p4143);
FA fa1663(ip_11_49,ip_12_48,ip_13_47,p4144,p4145);
FA fa1664(ip_14_46,ip_15_45,ip_16_44,p4146,p4147);
FA fa1665(ip_17_43,ip_18_42,ip_19_41,p4148,p4149);
FA fa1666(ip_20_40,ip_21_39,ip_22_38,p4150,p4151);
FA fa1667(ip_23_37,ip_24_36,ip_25_35,p4152,p4153);
HA ha409(ip_26_34,ip_27_33,p4154,p4155);
FA fa1668(ip_28_32,ip_29_31,ip_30_30,p4156,p4157);
FA fa1669(ip_31_29,ip_32_28,ip_33_27,p4158,p4159);
FA fa1670(ip_34_26,ip_35_25,ip_36_24,p4160,p4161);
HA ha410(ip_37_23,ip_38_22,p4162,p4163);
HA ha411(ip_39_21,ip_40_20,p4164,p4165);
HA ha412(ip_41_19,ip_42_18,p4166,p4167);
HA ha413(ip_43_17,ip_44_16,p4168,p4169);
FA fa1671(ip_45_15,ip_46_14,ip_47_13,p4170,p4171);
FA fa1672(ip_48_12,ip_49_11,ip_50_10,p4172,p4173);
FA fa1673(ip_51_9,ip_52_8,ip_53_7,p4174,p4175);
FA fa1674(ip_54_6,ip_55_5,ip_56_4,p4176,p4177);
HA ha414(ip_57_3,ip_58_2,p4178,p4179);
FA fa1675(ip_59_1,ip_60_0,p3990,p4180,p4181);
FA fa1676(p3998,p4012,p4022,p4182,p4183);
FA fa1677(p4024,p4141,p4155,p4184,p4185);
FA fa1678(p4163,p4165,p4167,p4186,p4187);
FA fa1679(p4169,p4179,p4030,p4188,p4189);
FA fa1680(p4034,p4137,p4139,p4190,p4191);
FA fa1681(p4143,p4145,p4147,p4192,p4193);
FA fa1682(p4149,p4151,p4153,p4194,p4195);
FA fa1683(p4157,p4159,p4161,p4196,p4197);
FA fa1684(p4171,p4173,p4175,p4198,p4199);
FA fa1685(p4177,p4181,p3986,p4200,p4201);
FA fa1686(p3988,p3992,p3994,p4202,p4203);
FA fa1687(p3996,p4000,p4002,p4204,p4205);
FA fa1688(p4004,p4006,p4008,p4206,p4207);
FA fa1689(p4010,p4014,p4016,p4208,p4209);
FA fa1690(p4018,p4020,p4026,p4210,p4211);
FA fa1691(p4028,p4183,p4185,p4212,p4213);
FA fa1692(p4187,p4189,p4032,p4214,p4215);
FA fa1693(p4036,p4052,p4056,p4216,p4217);
FA fa1694(p4191,p4193,p4195,p4218,p4219);
FA fa1695(p4197,p4199,p4201,p4220,p4221);
HA ha415(p4038,p4040,p4222,p4223);
FA fa1696(p4042,p4044,p4046,p4224,p4225);
FA fa1697(p4048,p4066,p4068,p4226,p4227);
FA fa1698(p4070,p4074,p4203,p4228,p4229);
FA fa1699(p4205,p4207,p4209,p4230,p4231);
FA fa1700(p4211,p4213,p4215,p4232,p4233);
FA fa1701(p4050,p4054,p4058,p4234,p4235);
FA fa1702(p4060,p4062,p4064,p4236,p4237);
FA fa1703(p4078,p4080,p4082,p4238,p4239);
FA fa1704(p4217,p4219,p4221,p4240,p4241);
FA fa1705(p4223,p4072,p4094,p4242,p4243);
FA fa1706(p4225,p4227,p4229,p4244,p4245);
HA ha416(p4231,p4233,p4246,p4247);
FA fa1707(p4076,p4084,p4086,p4248,p4249);
HA ha417(p4088,p4235,p4250,p4251);
FA fa1708(p4237,p4239,p4241,p4252,p4253);
FA fa1709(p4247,p4090,p4092,p4254,p4255);
FA fa1710(p4243,p4245,p4251,p4256,p4257);
FA fa1711(p4096,p4098,p4100,p4258,p4259);
HA ha418(p4102,p4249,p4260,p4261);
FA fa1712(p4253,p4104,p4106,p4262,p4263);
FA fa1713(p4255,p4257,p4261,p4264,p4265);
FA fa1714(p4108,p4110,p4259,p4266,p4267);
FA fa1715(p4112,p4114,p4263,p4268,p4269);
HA ha419(p4265,p4116,p4270,p4271);
FA fa1716(p4118,p4267,p4120,p4272,p4273);
FA fa1717(p4269,p4271,p4122,p4274,p4275);
FA fa1718(p4124,p4273,p4275,p4276,p4277);
FA fa1719(p4126,p4277,p4128,p4278,p4279);
FA fa1720(p4279,p4130,p4132,p4280,p4281);
FA fa1721(ip_0_61,ip_1_60,ip_2_59,p4282,p4283);
FA fa1722(ip_3_58,ip_4_57,ip_5_56,p4284,p4285);
FA fa1723(ip_6_55,ip_7_54,ip_8_53,p4286,p4287);
FA fa1724(ip_9_52,ip_10_51,ip_11_50,p4288,p4289);
FA fa1725(ip_12_49,ip_13_48,ip_14_47,p4290,p4291);
FA fa1726(ip_15_46,ip_16_45,ip_17_44,p4292,p4293);
FA fa1727(ip_18_43,ip_19_42,ip_20_41,p4294,p4295);
HA ha420(ip_21_40,ip_22_39,p4296,p4297);
FA fa1728(ip_23_38,ip_24_37,ip_25_36,p4298,p4299);
FA fa1729(ip_26_35,ip_27_34,ip_28_33,p4300,p4301);
FA fa1730(ip_29_32,ip_30_31,ip_31_30,p4302,p4303);
FA fa1731(ip_32_29,ip_33_28,ip_34_27,p4304,p4305);
FA fa1732(ip_35_26,ip_36_25,ip_37_24,p4306,p4307);
FA fa1733(ip_38_23,ip_39_22,ip_40_21,p4308,p4309);
FA fa1734(ip_41_20,ip_42_19,ip_43_18,p4310,p4311);
HA ha421(ip_44_17,ip_45_16,p4312,p4313);
FA fa1735(ip_46_15,ip_47_14,ip_48_13,p4314,p4315);
FA fa1736(ip_49_12,ip_50_11,ip_51_10,p4316,p4317);
FA fa1737(ip_52_9,ip_53_8,ip_54_7,p4318,p4319);
FA fa1738(ip_55_6,ip_56_5,ip_57_4,p4320,p4321);
FA fa1739(ip_58_3,ip_59_2,ip_60_1,p4322,p4323);
FA fa1740(ip_61_0,p4140,p4154,p4324,p4325);
FA fa1741(p4162,p4164,p4166,p4326,p4327);
FA fa1742(p4168,p4178,p4297,p4328,p4329);
HA ha422(p4313,p4283,p4330,p4331);
HA ha423(p4285,p4287,p4332,p4333);
FA fa1743(p4289,p4291,p4293,p4334,p4335);
FA fa1744(p4295,p4299,p4301,p4336,p4337);
FA fa1745(p4303,p4305,p4307,p4338,p4339);
FA fa1746(p4309,p4311,p4315,p4340,p4341);
FA fa1747(p4317,p4319,p4321,p4342,p4343);
FA fa1748(p4323,p4136,p4138,p4344,p4345);
FA fa1749(p4142,p4144,p4146,p4346,p4347);
FA fa1750(p4148,p4150,p4152,p4348,p4349);
FA fa1751(p4156,p4158,p4160,p4350,p4351);
FA fa1752(p4170,p4172,p4174,p4352,p4353);
HA ha424(p4176,p4180,p4354,p4355);
HA ha425(p4325,p4327,p4356,p4357);
HA ha426(p4329,p4331,p4358,p4359);
FA fa1753(p4333,p4182,p4184,p4360,p4361);
FA fa1754(p4186,p4188,p4335,p4362,p4363);
FA fa1755(p4337,p4339,p4341,p4364,p4365);
FA fa1756(p4343,p4355,p4357,p4366,p4367);
FA fa1757(p4359,p4190,p4192,p4368,p4369);
FA fa1758(p4194,p4196,p4198,p4370,p4371);
FA fa1759(p4200,p4345,p4347,p4372,p4373);
FA fa1760(p4349,p4351,p4353,p4374,p4375);
FA fa1761(p4202,p4204,p4206,p4376,p4377);
HA ha427(p4208,p4210,p4378,p4379);
HA ha428(p4212,p4214,p4380,p4381);
FA fa1762(p4222,p4361,p4363,p4382,p4383);
FA fa1763(p4365,p4367,p4216,p4384,p4385);
FA fa1764(p4218,p4220,p4369,p4386,p4387);
FA fa1765(p4371,p4373,p4375,p4388,p4389);
FA fa1766(p4379,p4381,p4224,p4390,p4391);
FA fa1767(p4226,p4228,p4230,p4392,p4393);
FA fa1768(p4232,p4246,p4377,p4394,p4395);
FA fa1769(p4383,p4385,p4234,p4396,p4397);
HA ha429(p4236,p4238,p4398,p4399);
FA fa1770(p4240,p4250,p4387,p4400,p4401);
FA fa1771(p4389,p4391,p4242,p4402,p4403);
HA ha430(p4244,p4393,p4404,p4405);
FA fa1772(p4395,p4397,p4399,p4406,p4407);
FA fa1773(p4248,p4252,p4260,p4408,p4409);
FA fa1774(p4401,p4403,p4405,p4410,p4411);
FA fa1775(p4254,p4256,p4407,p4412,p4413);
HA ha431(p4258,p4409,p4414,p4415);
FA fa1776(p4411,p4262,p4264,p4416,p4417);
FA fa1777(p4413,p4415,p4266,p4418,p4419);
FA fa1778(p4270,p4268,p4417,p4420,p4421);
FA fa1779(p4419,p4272,p4274,p4422,p4423);
FA fa1780(p4421,p4276,p4423,p4424,p4425);
FA fa1781(p4278,p4425,p4280,p4426,p4427);
FA fa1782(ip_0_62,ip_1_61,ip_2_60,p4428,p4429);
FA fa1783(ip_3_59,ip_4_58,ip_5_57,p4430,p4431);
FA fa1784(ip_6_56,ip_7_55,ip_8_54,p4432,p4433);
FA fa1785(ip_9_53,ip_10_52,ip_11_51,p4434,p4435);
FA fa1786(ip_12_50,ip_13_49,ip_14_48,p4436,p4437);
FA fa1787(ip_15_47,ip_16_46,ip_17_45,p4438,p4439);
FA fa1788(ip_18_44,ip_19_43,ip_20_42,p4440,p4441);
FA fa1789(ip_21_41,ip_22_40,ip_23_39,p4442,p4443);
FA fa1790(ip_24_38,ip_25_37,ip_26_36,p4444,p4445);
FA fa1791(ip_27_35,ip_28_34,ip_29_33,p4446,p4447);
HA ha432(ip_30_32,ip_31_31,p4448,p4449);
HA ha433(ip_32_30,ip_33_29,p4450,p4451);
FA fa1792(ip_34_28,ip_35_27,ip_36_26,p4452,p4453);
FA fa1793(ip_37_25,ip_38_24,ip_39_23,p4454,p4455);
HA ha434(ip_40_22,ip_41_21,p4456,p4457);
HA ha435(ip_42_20,ip_43_19,p4458,p4459);
FA fa1794(ip_44_18,ip_45_17,ip_46_16,p4460,p4461);
FA fa1795(ip_47_15,ip_48_14,ip_49_13,p4462,p4463);
FA fa1796(ip_50_12,ip_51_11,ip_52_10,p4464,p4465);
FA fa1797(ip_53_9,ip_54_8,ip_55_7,p4466,p4467);
FA fa1798(ip_56_6,ip_57_5,ip_58_4,p4468,p4469);
FA fa1799(ip_59_3,ip_60_2,ip_61_1,p4470,p4471);
FA fa1800(ip_62_0,p4296,p4312,p4472,p4473);
HA ha436(p4449,p4451,p4474,p4475);
HA ha437(p4457,p4459,p4476,p4477);
FA fa1801(p4429,p4431,p4433,p4478,p4479);
HA ha438(p4435,p4437,p4480,p4481);
FA fa1802(p4439,p4441,p4443,p4482,p4483);
FA fa1803(p4445,p4447,p4453,p4484,p4485);
FA fa1804(p4455,p4461,p4463,p4486,p4487);
FA fa1805(p4465,p4467,p4469,p4488,p4489);
FA fa1806(p4471,p4475,p4477,p4490,p4491);
FA fa1807(p4282,p4284,p4286,p4492,p4493);
FA fa1808(p4288,p4290,p4292,p4494,p4495);
HA ha439(p4294,p4298,p4496,p4497);
FA fa1809(p4300,p4302,p4304,p4498,p4499);
HA ha440(p4306,p4308,p4500,p4501);
FA fa1810(p4310,p4314,p4316,p4502,p4503);
FA fa1811(p4318,p4320,p4322,p4504,p4505);
FA fa1812(p4330,p4332,p4473,p4506,p4507);
FA fa1813(p4481,p4324,p4326,p4508,p4509);
FA fa1814(p4328,p4354,p4356,p4510,p4511);
FA fa1815(p4358,p4479,p4483,p4512,p4513);
FA fa1816(p4485,p4487,p4489,p4514,p4515);
FA fa1817(p4491,p4497,p4501,p4516,p4517);
HA ha441(p4334,p4336,p4518,p4519);
FA fa1818(p4338,p4340,p4342,p4520,p4521);
FA fa1819(p4493,p4495,p4499,p4522,p4523);
FA fa1820(p4503,p4505,p4507,p4524,p4525);
FA fa1821(p4344,p4346,p4348,p4526,p4527);
FA fa1822(p4350,p4352,p4509,p4528,p4529);
FA fa1823(p4511,p4513,p4515,p4530,p4531);
FA fa1824(p4517,p4519,p4360,p4532,p4533);
FA fa1825(p4362,p4364,p4366,p4534,p4535);
FA fa1826(p4378,p4380,p4521,p4536,p4537);
FA fa1827(p4523,p4525,p4368,p4538,p4539);
FA fa1828(p4370,p4372,p4374,p4540,p4541);
FA fa1829(p4527,p4529,p4531,p4542,p4543);
FA fa1830(p4533,p4376,p4382,p4544,p4545);
FA fa1831(p4384,p4535,p4537,p4546,p4547);
HA ha442(p4539,p4386,p4548,p4549);
HA ha443(p4388,p4390,p4550,p4551);
FA fa1832(p4398,p4541,p4543,p4552,p4553);
FA fa1833(p4392,p4394,p4396,p4554,p4555);
FA fa1834(p4404,p4545,p4547,p4556,p4557);
FA fa1835(p4549,p4551,p4400,p4558,p4559);
FA fa1836(p4402,p4553,p4406,p4560,p4561);
FA fa1837(p4555,p4557,p4559,p4562,p4563);
FA fa1838(p4408,p4410,p4414,p4564,p4565);
FA fa1839(p4561,p4412,p4563,p4566,p4567);
HA ha444(p4565,p4416,p4568,p4569);
FA fa1840(p4418,p4567,p4569,p4570,p4571);
FA fa1841(p4420,p4571,p4422,p4572,p4573);
FA fa1842(p4573,p4424,p4426,p4574,p4575);
FA fa1843(ip_0_63,ip_1_62,ip_2_61,p4576,p4577);
FA fa1844(ip_3_60,ip_4_59,ip_5_58,p4578,p4579);
FA fa1845(ip_6_57,ip_7_56,ip_8_55,p4580,p4581);
FA fa1846(ip_9_54,ip_10_53,ip_11_52,p4582,p4583);
FA fa1847(ip_12_51,ip_13_50,ip_14_49,p4584,p4585);
FA fa1848(ip_15_48,ip_16_47,ip_17_46,p4586,p4587);
FA fa1849(ip_18_45,ip_19_44,ip_20_43,p4588,p4589);
FA fa1850(ip_21_42,ip_22_41,ip_23_40,p4590,p4591);
FA fa1851(ip_24_39,ip_25_38,ip_26_37,p4592,p4593);
FA fa1852(ip_27_36,ip_28_35,ip_29_34,p4594,p4595);
FA fa1853(ip_30_33,ip_31_32,ip_32_31,p4596,p4597);
FA fa1854(ip_33_30,ip_34_29,ip_35_28,p4598,p4599);
FA fa1855(ip_36_27,ip_37_26,ip_38_25,p4600,p4601);
FA fa1856(ip_39_24,ip_40_23,ip_41_22,p4602,p4603);
FA fa1857(ip_42_21,ip_43_20,ip_44_19,p4604,p4605);
HA ha445(ip_45_18,ip_46_17,p4606,p4607);
FA fa1858(ip_47_16,ip_48_15,ip_49_14,p4608,p4609);
HA ha446(ip_50_13,ip_51_12,p4610,p4611);
FA fa1859(ip_52_11,ip_53_10,ip_54_9,p4612,p4613);
FA fa1860(ip_55_8,ip_56_7,ip_57_6,p4614,p4615);
HA ha447(ip_58_5,ip_59_4,p4616,p4617);
FA fa1861(ip_60_3,ip_61_2,ip_62_1,p4618,p4619);
HA ha448(ip_63_0,p4448,p4620,p4621);
FA fa1862(p4450,p4456,p4458,p4622,p4623);
HA ha449(p4607,p4611,p4624,p4625);
HA ha450(p4617,p4474,p4626,p4627);
FA fa1863(p4476,p4577,p4579,p4628,p4629);
FA fa1864(p4581,p4583,p4585,p4630,p4631);
FA fa1865(p4587,p4589,p4591,p4632,p4633);
HA ha451(p4593,p4595,p4634,p4635);
FA fa1866(p4597,p4599,p4601,p4636,p4637);
HA ha452(p4603,p4605,p4638,p4639);
FA fa1867(p4609,p4613,p4615,p4640,p4641);
FA fa1868(p4619,p4621,p4625,p4642,p4643);
FA fa1869(p4428,p4430,p4432,p4644,p4645);
FA fa1870(p4434,p4436,p4438,p4646,p4647);
HA ha453(p4440,p4442,p4648,p4649);
FA fa1871(p4444,p4446,p4452,p4650,p4651);
FA fa1872(p4454,p4460,p4462,p4652,p4653);
FA fa1873(p4464,p4466,p4468,p4654,p4655);
HA ha454(p4470,p4480,p4656,p4657);
HA ha455(p4623,p4627,p4658,p4659);
FA fa1874(p4635,p4639,p4472,p4660,p4661);
FA fa1875(p4496,p4500,p4629,p4662,p4663);
FA fa1876(p4631,p4633,p4637,p4664,p4665);
HA ha456(p4641,p4643,p4666,p4667);
FA fa1877(p4649,p4657,p4659,p4668,p4669);
FA fa1878(p4478,p4482,p4484,p4670,p4671);
FA fa1879(p4486,p4488,p4490,p4672,p4673);
FA fa1880(p4645,p4647,p4651,p4674,p4675);
FA fa1881(p4653,p4655,p4661,p4676,p4677);
FA fa1882(p4667,p4492,p4494,p4678,p4679);
HA ha457(p4498,p4502,p4680,p4681);
FA fa1883(p4504,p4506,p4518,p4682,p4683);
FA fa1884(p4663,p4665,p4669,p4684,p4685);
FA fa1885(p4508,p4510,p4512,p4686,p4687);
FA fa1886(p4514,p4516,p4671,p4688,p4689);
FA fa1887(p4673,p4675,p4677,p4690,p4691);
FA fa1888(p4681,p4520,p4522,p4692,p4693);
FA fa1889(p4524,p4679,p4683,p4694,p4695);
FA fa1890(p4685,p4526,p4528,p4696,p4697);
FA fa1891(p4530,p4532,p4687,p4698,p4699);
FA fa1892(p4689,p4691,p4534,p4700,p4701);
FA fa1893(p4536,p4538,p4693,p4702,p4703);
FA fa1894(p4695,p4540,p4542,p4704,p4705);
FA fa1895(p4548,p4550,p4697,p4706,p4707);
FA fa1896(p4699,p4701,p4544,p4708,p4709);
FA fa1897(p4546,p4703,p4552,p4710,p4711);
HA ha458(p4705,p4707,p4712,p4713);
HA ha459(p4709,p4554,p4714,p4715);
FA fa1898(p4556,p4558,p4711,p4716,p4717);
FA fa1899(p4713,p4560,p4715,p4718,p4719);
FA fa1900(p4562,p4717,p4564,p4720,p4721);
FA fa1901(p4719,p4566,p4568,p4722,p4723);
FA fa1902(p4721,p4570,p4723,p4724,p4725);
FA fa1903(p4572,p4725,p4574,p4726,p4727);
FA fa1904(ip_1_63,ip_2_62,ip_3_61,p4728,p4729);
FA fa1905(ip_4_60,ip_5_59,ip_6_58,p4730,p4731);
FA fa1906(ip_7_57,ip_8_56,ip_9_55,p4732,p4733);
FA fa1907(ip_10_54,ip_11_53,ip_12_52,p4734,p4735);
FA fa1908(ip_13_51,ip_14_50,ip_15_49,p4736,p4737);
FA fa1909(ip_16_48,ip_17_47,ip_18_46,p4738,p4739);
FA fa1910(ip_19_45,ip_20_44,ip_21_43,p4740,p4741);
FA fa1911(ip_22_42,ip_23_41,ip_24_40,p4742,p4743);
FA fa1912(ip_25_39,ip_26_38,ip_27_37,p4744,p4745);
FA fa1913(ip_28_36,ip_29_35,ip_30_34,p4746,p4747);
FA fa1914(ip_31_33,ip_32_32,ip_33_31,p4748,p4749);
HA ha460(ip_34_30,ip_35_29,p4750,p4751);
FA fa1915(ip_36_28,ip_37_27,ip_38_26,p4752,p4753);
FA fa1916(ip_39_25,ip_40_24,ip_41_23,p4754,p4755);
FA fa1917(ip_42_22,ip_43_21,ip_44_20,p4756,p4757);
FA fa1918(ip_45_19,ip_46_18,ip_47_17,p4758,p4759);
HA ha461(ip_48_16,ip_49_15,p4760,p4761);
FA fa1919(ip_50_14,ip_51_13,ip_52_12,p4762,p4763);
FA fa1920(ip_53_11,ip_54_10,ip_55_9,p4764,p4765);
FA fa1921(ip_56_8,ip_57_7,ip_58_6,p4766,p4767);
FA fa1922(ip_59_5,ip_60_4,ip_61_3,p4768,p4769);
FA fa1923(ip_62_2,ip_63_1,p4606,p4770,p4771);
HA ha462(p4610,p4616,p4772,p4773);
FA fa1924(p4751,p4761,p4620,p4774,p4775);
FA fa1925(p4624,p4729,p4731,p4776,p4777);
FA fa1926(p4733,p4735,p4737,p4778,p4779);
HA ha463(p4739,p4741,p4780,p4781);
FA fa1927(p4743,p4745,p4747,p4782,p4783);
HA ha464(p4749,p4753,p4784,p4785);
FA fa1928(p4755,p4757,p4759,p4786,p4787);
HA ha465(p4763,p4765,p4788,p4789);
HA ha466(p4767,p4769,p4790,p4791);
FA fa1929(p4771,p4773,p4576,p4792,p4793);
FA fa1930(p4578,p4580,p4582,p4794,p4795);
FA fa1931(p4584,p4586,p4588,p4796,p4797);
FA fa1932(p4590,p4592,p4594,p4798,p4799);
FA fa1933(p4596,p4598,p4600,p4800,p4801);
FA fa1934(p4602,p4604,p4608,p4802,p4803);
FA fa1935(p4612,p4614,p4618,p4804,p4805);
HA ha467(p4626,p4634,p4806,p4807);
FA fa1936(p4638,p4775,p4781,p4808,p4809);
HA ha468(p4785,p4789,p4810,p4811);
HA ha469(p4791,p4622,p4812,p4813);
FA fa1937(p4648,p4656,p4658,p4814,p4815);
HA ha470(p4777,p4779,p4816,p4817);
HA ha471(p4783,p4787,p4818,p4819);
HA ha472(p4793,p4807,p4820,p4821);
FA fa1938(p4811,p4628,p4630,p4822,p4823);
FA fa1939(p4632,p4636,p4640,p4824,p4825);
FA fa1940(p4642,p4666,p4795,p4826,p4827);
FA fa1941(p4797,p4799,p4801,p4828,p4829);
FA fa1942(p4803,p4805,p4809,p4830,p4831);
FA fa1943(p4813,p4817,p4819,p4832,p4833);
FA fa1944(p4821,p4644,p4646,p4834,p4835);
HA ha473(p4650,p4652,p4836,p4837);
FA fa1945(p4654,p4660,p4815,p4838,p4839);
HA ha474(p4662,p4664,p4840,p4841);
FA fa1946(p4668,p4680,p4823,p4842,p4843);
HA ha475(p4825,p4827,p4844,p4845);
FA fa1947(p4829,p4831,p4833,p4846,p4847);
FA fa1948(p4837,p4670,p4672,p4848,p4849);
FA fa1949(p4674,p4676,p4835,p4850,p4851);
FA fa1950(p4839,p4841,p4845,p4852,p4853);
FA fa1951(p4678,p4682,p4684,p4854,p4855);
FA fa1952(p4843,p4847,p4686,p4856,p4857);
FA fa1953(p4688,p4690,p4849,p4858,p4859);
HA ha476(p4851,p4853,p4860,p4861);
FA fa1954(p4692,p4694,p4855,p4862,p4863);
FA fa1955(p4857,p4861,p4696,p4864,p4865);
FA fa1956(p4698,p4700,p4859,p4866,p4867);
FA fa1957(p4702,p4863,p4865,p4868,p4869);
FA fa1958(p4704,p4706,p4708,p4870,p4871);
FA fa1959(p4712,p4867,p4710,p4872,p4873);
FA fa1960(p4714,p4869,p4871,p4874,p4875);
FA fa1961(p4873,p4716,p4875,p4876,p4877);
FA fa1962(p4718,p4720,p4877,p4878,p4879);
HA ha477(p4722,p4879,p4880,p4881);
FA fa1963(p4881,p4724,p4726,p4882,p4883);
HA ha478(ip_2_63,ip_3_62,p4884,p4885);
FA fa1964(ip_4_61,ip_5_60,ip_6_59,p4886,p4887);
FA fa1965(ip_7_58,ip_8_57,ip_9_56,p4888,p4889);
FA fa1966(ip_10_55,ip_11_54,ip_12_53,p4890,p4891);
HA ha479(ip_13_52,ip_14_51,p4892,p4893);
FA fa1967(ip_15_50,ip_16_49,ip_17_48,p4894,p4895);
FA fa1968(ip_18_47,ip_19_46,ip_20_45,p4896,p4897);
FA fa1969(ip_21_44,ip_22_43,ip_23_42,p4898,p4899);
FA fa1970(ip_24_41,ip_25_40,ip_26_39,p4900,p4901);
HA ha480(ip_27_38,ip_28_37,p4902,p4903);
FA fa1971(ip_29_36,ip_30_35,ip_31_34,p4904,p4905);
FA fa1972(ip_32_33,ip_33_32,ip_34_31,p4906,p4907);
FA fa1973(ip_35_30,ip_36_29,ip_37_28,p4908,p4909);
FA fa1974(ip_38_27,ip_39_26,ip_40_25,p4910,p4911);
FA fa1975(ip_41_24,ip_42_23,ip_43_22,p4912,p4913);
FA fa1976(ip_44_21,ip_45_20,ip_46_19,p4914,p4915);
HA ha481(ip_47_18,ip_48_17,p4916,p4917);
FA fa1977(ip_49_16,ip_50_15,ip_51_14,p4918,p4919);
FA fa1978(ip_52_13,ip_53_12,ip_54_11,p4920,p4921);
FA fa1979(ip_55_10,ip_56_9,ip_57_8,p4922,p4923);
FA fa1980(ip_58_7,ip_59_6,ip_60_5,p4924,p4925);
FA fa1981(ip_61_4,ip_62_3,ip_63_2,p4926,p4927);
FA fa1982(p4750,p4760,p4885,p4928,p4929);
FA fa1983(p4893,p4903,p4917,p4930,p4931);
HA ha482(p4772,p4887,p4932,p4933);
FA fa1984(p4889,p4891,p4895,p4934,p4935);
HA ha483(p4897,p4899,p4936,p4937);
HA ha484(p4901,p4905,p4938,p4939);
FA fa1985(p4907,p4909,p4911,p4940,p4941);
FA fa1986(p4913,p4915,p4919,p4942,p4943);
FA fa1987(p4921,p4923,p4925,p4944,p4945);
HA ha485(p4927,p4728,p4946,p4947);
FA fa1988(p4730,p4732,p4734,p4948,p4949);
FA fa1989(p4736,p4738,p4740,p4950,p4951);
FA fa1990(p4742,p4744,p4746,p4952,p4953);
FA fa1991(p4748,p4752,p4754,p4954,p4955);
FA fa1992(p4756,p4758,p4762,p4956,p4957);
FA fa1993(p4764,p4766,p4768,p4958,p4959);
FA fa1994(p4770,p4780,p4784,p4960,p4961);
FA fa1995(p4788,p4790,p4929,p4962,p4963);
FA fa1996(p4931,p4933,p4937,p4964,p4965);
HA ha486(p4939,p4774,p4966,p4967);
FA fa1997(p4806,p4810,p4935,p4968,p4969);
FA fa1998(p4941,p4943,p4945,p4970,p4971);
FA fa1999(p4947,p4776,p4778,p4972,p4973);
FA fa2000(p4782,p4786,p4792,p4974,p4975);
FA fa2001(p4812,p4816,p4818,p4976,p4977);
FA fa2002(p4820,p4949,p4951,p4978,p4979);
FA fa2003(p4953,p4955,p4957,p4980,p4981);
FA fa2004(p4959,p4961,p4963,p4982,p4983);
HA ha487(p4965,p4967,p4984,p4985);
FA fa2005(p4794,p4796,p4798,p4986,p4987);
FA fa2006(p4800,p4802,p4804,p4988,p4989);
FA fa2007(p4808,p4969,p4971,p4990,p4991);
FA fa2008(p4985,p4814,p4836,p4992,p4993);
FA fa2009(p4973,p4975,p4977,p4994,p4995);
FA fa2010(p4979,p4981,p4983,p4996,p4997);
FA fa2011(p4822,p4824,p4826,p4998,p4999);
FA fa2012(p4828,p4830,p4832,p5000,p5001);
FA fa2013(p4840,p4844,p4987,p5002,p5003);
HA ha488(p4989,p4991,p5004,p5005);
FA fa2014(p4834,p4838,p4993,p5006,p5007);
HA ha489(p4995,p4997,p5008,p5009);
FA fa2015(p5005,p4842,p4846,p5010,p5011);
HA ha490(p4999,p5001,p5012,p5013);
FA fa2016(p5003,p5009,p4848,p5014,p5015);
FA fa2017(p4850,p4852,p4860,p5016,p5017);
HA ha491(p5007,p5013,p5018,p5019);
FA fa2018(p4854,p4856,p5011,p5020,p5021);
FA fa2019(p5015,p5019,p4858,p5022,p5023);
HA ha492(p5017,p4862,p5024,p5025);
FA fa2020(p4864,p5021,p5023,p5026,p5027);
FA fa2021(p4866,p5025,p4868,p5028,p5029);
FA fa2022(p5027,p4870,p4872,p5030,p5031);
FA fa2023(p5029,p4874,p5031,p5032,p5033);
FA fa2024(p4876,p5033,p4878,p5034,p5035);
FA fa2025(p4880,p5035,p4882,p5036,p5037);
HA ha493(ip_3_63,ip_4_62,p5038,p5039);
FA fa2026(ip_5_61,ip_6_60,ip_7_59,p5040,p5041);
FA fa2027(ip_8_58,ip_9_57,ip_10_56,p5042,p5043);
FA fa2028(ip_11_55,ip_12_54,ip_13_53,p5044,p5045);
FA fa2029(ip_14_52,ip_15_51,ip_16_50,p5046,p5047);
FA fa2030(ip_17_49,ip_18_48,ip_19_47,p5048,p5049);
FA fa2031(ip_20_46,ip_21_45,ip_22_44,p5050,p5051);
FA fa2032(ip_23_43,ip_24_42,ip_25_41,p5052,p5053);
FA fa2033(ip_26_40,ip_27_39,ip_28_38,p5054,p5055);
HA ha494(ip_29_37,ip_30_36,p5056,p5057);
FA fa2034(ip_31_35,ip_32_34,ip_33_33,p5058,p5059);
FA fa2035(ip_34_32,ip_35_31,ip_36_30,p5060,p5061);
FA fa2036(ip_37_29,ip_38_28,ip_39_27,p5062,p5063);
FA fa2037(ip_40_26,ip_41_25,ip_42_24,p5064,p5065);
FA fa2038(ip_43_23,ip_44_22,ip_45_21,p5066,p5067);
FA fa2039(ip_46_20,ip_47_19,ip_48_18,p5068,p5069);
FA fa2040(ip_49_17,ip_50_16,ip_51_15,p5070,p5071);
FA fa2041(ip_52_14,ip_53_13,ip_54_12,p5072,p5073);
FA fa2042(ip_55_11,ip_56_10,ip_57_9,p5074,p5075);
FA fa2043(ip_58_8,ip_59_7,ip_60_6,p5076,p5077);
HA ha495(ip_61_5,ip_62_4,p5078,p5079);
FA fa2044(ip_63_3,p4884,p4892,p5080,p5081);
HA ha496(p4902,p4916,p5082,p5083);
HA ha497(p5039,p5057,p5084,p5085);
FA fa2045(p5079,p5041,p5043,p5086,p5087);
FA fa2046(p5045,p5047,p5049,p5088,p5089);
FA fa2047(p5051,p5053,p5055,p5090,p5091);
FA fa2048(p5059,p5061,p5063,p5092,p5093);
FA fa2049(p5065,p5067,p5069,p5094,p5095);
FA fa2050(p5071,p5073,p5075,p5096,p5097);
HA ha498(p5077,p5083,p5098,p5099);
FA fa2051(p5085,p4886,p4888,p5100,p5101);
HA ha499(p4890,p4894,p5102,p5103);
HA ha500(p4896,p4898,p5104,p5105);
FA fa2052(p4900,p4904,p4906,p5106,p5107);
FA fa2053(p4908,p4910,p4912,p5108,p5109);
FA fa2054(p4914,p4918,p4920,p5110,p5111);
FA fa2055(p4922,p4924,p4926,p5112,p5113);
FA fa2056(p4932,p4936,p4938,p5114,p5115);
HA ha501(p5081,p5099,p5116,p5117);
FA fa2057(p4928,p4930,p4946,p5118,p5119);
FA fa2058(p5087,p5089,p5091,p5120,p5121);
HA ha502(p5093,p5095,p5122,p5123);
FA fa2059(p5097,p5103,p5105,p5124,p5125);
HA ha503(p5117,p4934,p5126,p5127);
HA ha504(p4940,p4942,p5128,p5129);
FA fa2060(p4944,p4966,p5101,p5130,p5131);
FA fa2061(p5107,p5109,p5111,p5132,p5133);
FA fa2062(p5113,p5115,p5123,p5134,p5135);
FA fa2063(p4948,p4950,p4952,p5136,p5137);
FA fa2064(p4954,p4956,p4958,p5138,p5139);
HA ha505(p4960,p4962,p5140,p5141);
FA fa2065(p4964,p4984,p5119,p5142,p5143);
HA ha506(p5121,p5125,p5144,p5145);
FA fa2066(p5127,p5129,p4968,p5146,p5147);
FA fa2067(p4970,p5131,p5133,p5148,p5149);
FA fa2068(p5135,p5141,p5145,p5150,p5151);
HA ha507(p4972,p4974,p5152,p5153);
FA fa2069(p4976,p4978,p4980,p5154,p5155);
FA fa2070(p4982,p5137,p5139,p5156,p5157);
FA fa2071(p5143,p5147,p4986,p5158,p5159);
HA ha508(p4988,p4990,p5160,p5161);
FA fa2072(p5004,p5149,p5151,p5162,p5163);
FA fa2073(p5153,p4992,p4994,p5164,p5165);
FA fa2074(p4996,p5008,p5155,p5166,p5167);
FA fa2075(p5157,p5159,p5161,p5168,p5169);
HA ha509(p4998,p5000,p5170,p5171);
FA fa2076(p5002,p5012,p5163,p5172,p5173);
FA fa2077(p5006,p5018,p5165,p5174,p5175);
FA fa2078(p5167,p5169,p5171,p5176,p5177);
FA fa2079(p5010,p5014,p5173,p5178,p5179);
FA fa2080(p5016,p5175,p5177,p5180,p5181);
FA fa2081(p5020,p5022,p5024,p5182,p5183);
HA ha510(p5179,p5181,p5184,p5185);
FA fa2082(p5026,p5183,p5185,p5186,p5187);
FA fa2083(p5028,p5187,p5030,p5188,p5189);
FA fa2084(p5032,p5189,p5034,p5190,p5191);
FA fa2085(ip_4_63,ip_5_62,ip_6_61,p5192,p5193);
FA fa2086(ip_7_60,ip_8_59,ip_9_58,p5194,p5195);
HA ha511(ip_10_57,ip_11_56,p5196,p5197);
HA ha512(ip_12_55,ip_13_54,p5198,p5199);
HA ha513(ip_14_53,ip_15_52,p5200,p5201);
FA fa2087(ip_16_51,ip_17_50,ip_18_49,p5202,p5203);
HA ha514(ip_19_48,ip_20_47,p5204,p5205);
FA fa2088(ip_21_46,ip_22_45,ip_23_44,p5206,p5207);
FA fa2089(ip_24_43,ip_25_42,ip_26_41,p5208,p5209);
FA fa2090(ip_27_40,ip_28_39,ip_29_38,p5210,p5211);
HA ha515(ip_30_37,ip_31_36,p5212,p5213);
FA fa2091(ip_32_35,ip_33_34,ip_34_33,p5214,p5215);
HA ha516(ip_35_32,ip_36_31,p5216,p5217);
FA fa2092(ip_37_30,ip_38_29,ip_39_28,p5218,p5219);
FA fa2093(ip_40_27,ip_41_26,ip_42_25,p5220,p5221);
FA fa2094(ip_43_24,ip_44_23,ip_45_22,p5222,p5223);
FA fa2095(ip_46_21,ip_47_20,ip_48_19,p5224,p5225);
FA fa2096(ip_49_18,ip_50_17,ip_51_16,p5226,p5227);
HA ha517(ip_52_15,ip_53_14,p5228,p5229);
HA ha518(ip_54_13,ip_55_12,p5230,p5231);
FA fa2097(ip_56_11,ip_57_10,ip_58_9,p5232,p5233);
FA fa2098(ip_59_8,ip_60_7,ip_61_6,p5234,p5235);
FA fa2099(ip_62_5,ip_63_4,p5038,p5236,p5237);
FA fa2100(p5056,p5078,p5197,p5238,p5239);
FA fa2101(p5199,p5201,p5205,p5240,p5241);
HA ha519(p5213,p5217,p5242,p5243);
FA fa2102(p5229,p5231,p5082,p5244,p5245);
FA fa2103(p5084,p5193,p5195,p5246,p5247);
FA fa2104(p5203,p5207,p5209,p5248,p5249);
FA fa2105(p5211,p5215,p5219,p5250,p5251);
HA ha520(p5221,p5223,p5252,p5253);
HA ha521(p5225,p5227,p5254,p5255);
HA ha522(p5233,p5235,p5256,p5257);
FA fa2106(p5237,p5243,p5040,p5258,p5259);
FA fa2107(p5042,p5044,p5046,p5260,p5261);
HA ha523(p5048,p5050,p5262,p5263);
FA fa2108(p5052,p5054,p5058,p5264,p5265);
FA fa2109(p5060,p5062,p5064,p5266,p5267);
FA fa2110(p5066,p5068,p5070,p5268,p5269);
FA fa2111(p5072,p5074,p5076,p5270,p5271);
FA fa2112(p5098,p5239,p5241,p5272,p5273);
FA fa2113(p5245,p5253,p5255,p5274,p5275);
HA ha524(p5257,p5080,p5276,p5277);
FA fa2114(p5102,p5104,p5116,p5278,p5279);
FA fa2115(p5247,p5249,p5251,p5280,p5281);
FA fa2116(p5259,p5263,p5086,p5282,p5283);
FA fa2117(p5088,p5090,p5092,p5284,p5285);
HA ha525(p5094,p5096,p5286,p5287);
HA ha526(p5122,p5261,p5288,p5289);
FA fa2118(p5265,p5267,p5269,p5290,p5291);
HA ha527(p5271,p5273,p5292,p5293);
FA fa2119(p5275,p5277,p5100,p5294,p5295);
FA fa2120(p5106,p5108,p5110,p5296,p5297);
FA fa2121(p5112,p5114,p5126,p5298,p5299);
FA fa2122(p5128,p5279,p5281,p5300,p5301);
FA fa2123(p5283,p5287,p5289,p5302,p5303);
FA fa2124(p5293,p5118,p5120,p5304,p5305);
FA fa2125(p5124,p5140,p5144,p5306,p5307);
FA fa2126(p5285,p5291,p5295,p5308,p5309);
HA ha528(p5130,p5132,p5310,p5311);
FA fa2127(p5134,p5297,p5299,p5312,p5313);
FA fa2128(p5301,p5303,p5136,p5314,p5315);
FA fa2129(p5138,p5142,p5146,p5316,p5317);
FA fa2130(p5152,p5305,p5307,p5318,p5319);
FA fa2131(p5309,p5311,p5148,p5320,p5321);
HA ha529(p5150,p5160,p5322,p5323);
FA fa2132(p5313,p5315,p5154,p5324,p5325);
FA fa2133(p5156,p5158,p5317,p5326,p5327);
FA fa2134(p5319,p5321,p5323,p5328,p5329);
FA fa2135(p5162,p5170,p5325,p5330,p5331);
FA fa2136(p5164,p5166,p5168,p5332,p5333);
FA fa2137(p5327,p5329,p5172,p5334,p5335);
FA fa2138(p5331,p5174,p5176,p5336,p5337);
FA fa2139(p5333,p5335,p5178,p5338,p5339);
FA fa2140(p5180,p5184,p5337,p5340,p5341);
FA fa2141(p5339,p5182,p5341,p5342,p5343);
FA fa2142(p5186,p5343,p5188,p5344,p5345);
HA ha530(ip_5_63,ip_6_62,p5346,p5347);
HA ha531(ip_7_61,ip_8_60,p5348,p5349);
FA fa2143(ip_9_59,ip_10_58,ip_11_57,p5350,p5351);
HA ha532(ip_12_56,ip_13_55,p5352,p5353);
FA fa2144(ip_14_54,ip_15_53,ip_16_52,p5354,p5355);
FA fa2145(ip_17_51,ip_18_50,ip_19_49,p5356,p5357);
FA fa2146(ip_20_48,ip_21_47,ip_22_46,p5358,p5359);
HA ha533(ip_23_45,ip_24_44,p5360,p5361);
FA fa2147(ip_25_43,ip_26_42,ip_27_41,p5362,p5363);
FA fa2148(ip_28_40,ip_29_39,ip_30_38,p5364,p5365);
FA fa2149(ip_31_37,ip_32_36,ip_33_35,p5366,p5367);
FA fa2150(ip_34_34,ip_35_33,ip_36_32,p5368,p5369);
FA fa2151(ip_37_31,ip_38_30,ip_39_29,p5370,p5371);
FA fa2152(ip_40_28,ip_41_27,ip_42_26,p5372,p5373);
FA fa2153(ip_43_25,ip_44_24,ip_45_23,p5374,p5375);
FA fa2154(ip_46_22,ip_47_21,ip_48_20,p5376,p5377);
FA fa2155(ip_49_19,ip_50_18,ip_51_17,p5378,p5379);
FA fa2156(ip_52_16,ip_53_15,ip_54_14,p5380,p5381);
HA ha534(ip_55_13,ip_56_12,p5382,p5383);
FA fa2157(ip_57_11,ip_58_10,ip_59_9,p5384,p5385);
FA fa2158(ip_60_8,ip_61_7,ip_62_6,p5386,p5387);
FA fa2159(ip_63_5,p5196,p5198,p5388,p5389);
FA fa2160(p5200,p5204,p5212,p5390,p5391);
FA fa2161(p5216,p5228,p5230,p5392,p5393);
FA fa2162(p5347,p5349,p5353,p5394,p5395);
FA fa2163(p5361,p5383,p5242,p5396,p5397);
FA fa2164(p5351,p5355,p5357,p5398,p5399);
FA fa2165(p5359,p5363,p5365,p5400,p5401);
FA fa2166(p5367,p5369,p5371,p5402,p5403);
FA fa2167(p5373,p5375,p5377,p5404,p5405);
FA fa2168(p5379,p5381,p5385,p5406,p5407);
FA fa2169(p5387,p5192,p5194,p5408,p5409);
FA fa2170(p5202,p5206,p5208,p5410,p5411);
FA fa2171(p5210,p5214,p5218,p5412,p5413);
HA ha535(p5220,p5222,p5414,p5415);
FA fa2172(p5224,p5226,p5232,p5416,p5417);
HA ha536(p5234,p5236,p5418,p5419);
FA fa2173(p5252,p5254,p5256,p5420,p5421);
HA ha537(p5389,p5391,p5422,p5423);
FA fa2174(p5393,p5395,p5397,p5424,p5425);
FA fa2175(p5238,p5240,p5244,p5426,p5427);
FA fa2176(p5262,p5399,p5401,p5428,p5429);
FA fa2177(p5403,p5405,p5407,p5430,p5431);
FA fa2178(p5415,p5419,p5423,p5432,p5433);
HA ha538(p5246,p5248,p5434,p5435);
HA ha539(p5250,p5258,p5436,p5437);
FA fa2179(p5276,p5409,p5411,p5438,p5439);
FA fa2180(p5413,p5417,p5421,p5440,p5441);
FA fa2181(p5425,p5260,p5264,p5442,p5443);
FA fa2182(p5266,p5268,p5270,p5444,p5445);
HA ha540(p5272,p5274,p5446,p5447);
FA fa2183(p5286,p5288,p5292,p5448,p5449);
FA fa2184(p5427,p5429,p5431,p5450,p5451);
FA fa2185(p5433,p5435,p5437,p5452,p5453);
FA fa2186(p5278,p5280,p5282,p5454,p5455);
FA fa2187(p5439,p5441,p5447,p5456,p5457);
FA fa2188(p5284,p5290,p5294,p5458,p5459);
HA ha541(p5443,p5445,p5460,p5461);
FA fa2189(p5449,p5451,p5453,p5462,p5463);
FA fa2190(p5296,p5298,p5300,p5464,p5465);
FA fa2191(p5302,p5310,p5455,p5466,p5467);
FA fa2192(p5457,p5461,p5304,p5468,p5469);
FA fa2193(p5306,p5308,p5459,p5470,p5471);
FA fa2194(p5463,p5312,p5314,p5472,p5473);
FA fa2195(p5322,p5465,p5467,p5474,p5475);
FA fa2196(p5469,p5316,p5318,p5476,p5477);
FA fa2197(p5320,p5471,p5324,p5478,p5479);
FA fa2198(p5473,p5475,p5326,p5480,p5481);
FA fa2199(p5328,p5477,p5479,p5482,p5483);
FA fa2200(p5330,p5481,p5332,p5484,p5485);
HA ha542(p5334,p5483,p5486,p5487);
FA fa2201(p5485,p5487,p5336,p5488,p5489);
HA ha543(p5338,p5489,p5490,p5491);
FA fa2202(p5340,p5491,p5342,p5492,p5493);
HA ha544(ip_6_63,ip_7_62,p5494,p5495);
FA fa2203(ip_8_61,ip_9_60,ip_10_59,p5496,p5497);
FA fa2204(ip_11_58,ip_12_57,ip_13_56,p5498,p5499);
FA fa2205(ip_14_55,ip_15_54,ip_16_53,p5500,p5501);
HA ha545(ip_17_52,ip_18_51,p5502,p5503);
HA ha546(ip_19_50,ip_20_49,p5504,p5505);
FA fa2206(ip_21_48,ip_22_47,ip_23_46,p5506,p5507);
FA fa2207(ip_24_45,ip_25_44,ip_26_43,p5508,p5509);
HA ha547(ip_27_42,ip_28_41,p5510,p5511);
HA ha548(ip_29_40,ip_30_39,p5512,p5513);
FA fa2208(ip_31_38,ip_32_37,ip_33_36,p5514,p5515);
FA fa2209(ip_34_35,ip_35_34,ip_36_33,p5516,p5517);
FA fa2210(ip_37_32,ip_38_31,ip_39_30,p5518,p5519);
FA fa2211(ip_40_29,ip_41_28,ip_42_27,p5520,p5521);
FA fa2212(ip_43_26,ip_44_25,ip_45_24,p5522,p5523);
FA fa2213(ip_46_23,ip_47_22,ip_48_21,p5524,p5525);
HA ha549(ip_49_20,ip_50_19,p5526,p5527);
FA fa2214(ip_51_18,ip_52_17,ip_53_16,p5528,p5529);
FA fa2215(ip_54_15,ip_55_14,ip_56_13,p5530,p5531);
FA fa2216(ip_57_12,ip_58_11,ip_59_10,p5532,p5533);
FA fa2217(ip_60_9,ip_61_8,ip_62_7,p5534,p5535);
FA fa2218(ip_63_6,p5346,p5348,p5536,p5537);
FA fa2219(p5352,p5360,p5382,p5538,p5539);
HA ha550(p5495,p5503,p5540,p5541);
FA fa2220(p5505,p5511,p5513,p5542,p5543);
FA fa2221(p5527,p5497,p5499,p5544,p5545);
HA ha551(p5501,p5507,p5546,p5547);
HA ha552(p5509,p5515,p5548,p5549);
FA fa2222(p5517,p5519,p5521,p5550,p5551);
FA fa2223(p5523,p5525,p5529,p5552,p5553);
FA fa2224(p5531,p5533,p5535,p5554,p5555);
FA fa2225(p5541,p5350,p5354,p5556,p5557);
FA fa2226(p5356,p5358,p5362,p5558,p5559);
HA ha553(p5364,p5366,p5560,p5561);
FA fa2227(p5368,p5370,p5372,p5562,p5563);
FA fa2228(p5374,p5376,p5378,p5564,p5565);
FA fa2229(p5380,p5384,p5386,p5566,p5567);
FA fa2230(p5537,p5539,p5543,p5568,p5569);
FA fa2231(p5547,p5549,p5388,p5570,p5571);
FA fa2232(p5390,p5392,p5394,p5572,p5573);
FA fa2233(p5396,p5414,p5418,p5574,p5575);
HA ha554(p5422,p5545,p5576,p5577);
FA fa2234(p5551,p5553,p5555,p5578,p5579);
FA fa2235(p5561,p5398,p5400,p5580,p5581);
FA fa2236(p5402,p5404,p5406,p5582,p5583);
FA fa2237(p5557,p5559,p5563,p5584,p5585);
HA ha555(p5565,p5567,p5586,p5587);
FA fa2238(p5569,p5571,p5577,p5588,p5589);
FA fa2239(p5408,p5410,p5412,p5590,p5591);
FA fa2240(p5416,p5420,p5424,p5592,p5593);
FA fa2241(p5434,p5436,p5573,p5594,p5595);
FA fa2242(p5575,p5579,p5587,p5596,p5597);
FA fa2243(p5426,p5428,p5430,p5598,p5599);
FA fa2244(p5432,p5446,p5581,p5600,p5601);
FA fa2245(p5583,p5585,p5589,p5602,p5603);
FA fa2246(p5438,p5440,p5591,p5604,p5605);
HA ha556(p5593,p5595,p5606,p5607);
HA ha557(p5597,p5442,p5608,p5609);
FA fa2247(p5444,p5448,p5450,p5610,p5611);
HA ha558(p5452,p5460,p5612,p5613);
FA fa2248(p5599,p5601,p5603,p5614,p5615);
FA fa2249(p5607,p5454,p5456,p5616,p5617);
HA ha559(p5605,p5609,p5618,p5619);
FA fa2250(p5613,p5458,p5462,p5620,p5621);
FA fa2251(p5611,p5615,p5619,p5622,p5623);
FA fa2252(p5464,p5466,p5468,p5624,p5625);
FA fa2253(p5617,p5470,p5621,p5626,p5627);
FA fa2254(p5623,p5472,p5474,p5628,p5629);
FA fa2255(p5625,p5476,p5478,p5630,p5631);
FA fa2256(p5627,p5480,p5629,p5632,p5633);
FA fa2257(p5482,p5486,p5631,p5634,p5635);
FA fa2258(p5484,p5633,p5635,p5636,p5637);
HA ha560(p5488,p5490,p5638,p5639);
FA fa2259(p5637,p5639,p5492,p5640,p5641);
HA ha561(ip_7_63,ip_8_62,p5642,p5643);
HA ha562(ip_9_61,ip_10_60,p5644,p5645);
FA fa2260(ip_11_59,ip_12_58,ip_13_57,p5646,p5647);
FA fa2261(ip_14_56,ip_15_55,ip_16_54,p5648,p5649);
FA fa2262(ip_17_53,ip_18_52,ip_19_51,p5650,p5651);
FA fa2263(ip_20_50,ip_21_49,ip_22_48,p5652,p5653);
FA fa2264(ip_23_47,ip_24_46,ip_25_45,p5654,p5655);
FA fa2265(ip_26_44,ip_27_43,ip_28_42,p5656,p5657);
FA fa2266(ip_29_41,ip_30_40,ip_31_39,p5658,p5659);
HA ha563(ip_32_38,ip_33_37,p5660,p5661);
FA fa2267(ip_34_36,ip_35_35,ip_36_34,p5662,p5663);
FA fa2268(ip_37_33,ip_38_32,ip_39_31,p5664,p5665);
FA fa2269(ip_40_30,ip_41_29,ip_42_28,p5666,p5667);
FA fa2270(ip_43_27,ip_44_26,ip_45_25,p5668,p5669);
HA ha564(ip_46_24,ip_47_23,p5670,p5671);
HA ha565(ip_48_22,ip_49_21,p5672,p5673);
FA fa2271(ip_50_20,ip_51_19,ip_52_18,p5674,p5675);
FA fa2272(ip_53_17,ip_54_16,ip_55_15,p5676,p5677);
HA ha566(ip_56_14,ip_57_13,p5678,p5679);
FA fa2273(ip_58_12,ip_59_11,ip_60_10,p5680,p5681);
FA fa2274(ip_61_9,ip_62_8,ip_63_7,p5682,p5683);
FA fa2275(p5494,p5502,p5504,p5684,p5685);
HA ha567(p5510,p5512,p5686,p5687);
FA fa2276(p5526,p5643,p5645,p5688,p5689);
FA fa2277(p5661,p5671,p5673,p5690,p5691);
FA fa2278(p5679,p5540,p5647,p5692,p5693);
FA fa2279(p5649,p5651,p5653,p5694,p5695);
HA ha568(p5655,p5657,p5696,p5697);
HA ha569(p5659,p5663,p5698,p5699);
FA fa2280(p5665,p5667,p5669,p5700,p5701);
HA ha570(p5675,p5677,p5702,p5703);
HA ha571(p5681,p5683,p5704,p5705);
FA fa2281(p5687,p5496,p5498,p5706,p5707);
HA ha572(p5500,p5506,p5708,p5709);
FA fa2282(p5508,p5514,p5516,p5710,p5711);
FA fa2283(p5518,p5520,p5522,p5712,p5713);
FA fa2284(p5524,p5528,p5530,p5714,p5715);
HA ha573(p5532,p5534,p5716,p5717);
HA ha574(p5546,p5548,p5718,p5719);
HA ha575(p5685,p5689,p5720,p5721);
HA ha576(p5691,p5697,p5722,p5723);
FA fa2285(p5699,p5703,p5705,p5724,p5725);
FA fa2286(p5536,p5538,p5542,p5726,p5727);
HA ha577(p5560,p5693,p5728,p5729);
FA fa2287(p5695,p5701,p5709,p5730,p5731);
FA fa2288(p5717,p5719,p5721,p5732,p5733);
HA ha578(p5723,p5544,p5734,p5735);
HA ha579(p5550,p5552,p5736,p5737);
FA fa2289(p5554,p5576,p5707,p5738,p5739);
FA fa2290(p5711,p5713,p5715,p5740,p5741);
FA fa2291(p5725,p5729,p5556,p5742,p5743);
FA fa2292(p5558,p5562,p5564,p5744,p5745);
FA fa2293(p5566,p5568,p5570,p5746,p5747);
HA ha580(p5586,p5727,p5748,p5749);
HA ha581(p5731,p5733,p5750,p5751);
FA fa2294(p5735,p5737,p5572,p5752,p5753);
FA fa2295(p5574,p5578,p5739,p5754,p5755);
FA fa2296(p5741,p5743,p5749,p5756,p5757);
FA fa2297(p5751,p5580,p5582,p5758,p5759);
FA fa2298(p5584,p5588,p5745,p5760,p5761);
FA fa2299(p5747,p5753,p5590,p5762,p5763);
FA fa2300(p5592,p5594,p5596,p5764,p5765);
FA fa2301(p5606,p5755,p5757,p5766,p5767);
FA fa2302(p5598,p5600,p5602,p5768,p5769);
FA fa2303(p5608,p5612,p5759,p5770,p5771);
HA ha582(p5761,p5763,p5772,p5773);
FA fa2304(p5604,p5618,p5765,p5774,p5775);
FA fa2305(p5767,p5773,p5610,p5776,p5777);
FA fa2306(p5614,p5769,p5771,p5778,p5779);
HA ha583(p5616,p5775,p5780,p5781);
FA fa2307(p5777,p5620,p5622,p5782,p5783);
FA fa2308(p5779,p5781,p5624,p5784,p5785);
FA fa2309(p5626,p5783,p5785,p5786,p5787);
HA ha584(p5628,p5630,p5788,p5789);
HA ha585(p5787,p5632,p5790,p5791);
FA fa2310(p5789,p5634,p5791,p5792,p5793);
HA ha586(p5636,p5638,p5794,p5795);
FA fa2311(p5793,p5795,p5640,p5796,p5797);
FA fa2312(ip_8_63,ip_9_62,ip_10_61,p5798,p5799);
FA fa2313(ip_11_60,ip_12_59,ip_13_58,p5800,p5801);
FA fa2314(ip_14_57,ip_15_56,ip_16_55,p5802,p5803);
FA fa2315(ip_17_54,ip_18_53,ip_19_52,p5804,p5805);
FA fa2316(ip_20_51,ip_21_50,ip_22_49,p5806,p5807);
FA fa2317(ip_23_48,ip_24_47,ip_25_46,p5808,p5809);
FA fa2318(ip_26_45,ip_27_44,ip_28_43,p5810,p5811);
FA fa2319(ip_29_42,ip_30_41,ip_31_40,p5812,p5813);
FA fa2320(ip_32_39,ip_33_38,ip_34_37,p5814,p5815);
FA fa2321(ip_35_36,ip_36_35,ip_37_34,p5816,p5817);
FA fa2322(ip_38_33,ip_39_32,ip_40_31,p5818,p5819);
FA fa2323(ip_41_30,ip_42_29,ip_43_28,p5820,p5821);
FA fa2324(ip_44_27,ip_45_26,ip_46_25,p5822,p5823);
FA fa2325(ip_47_24,ip_48_23,ip_49_22,p5824,p5825);
HA ha587(ip_50_21,ip_51_20,p5826,p5827);
FA fa2326(ip_52_19,ip_53_18,ip_54_17,p5828,p5829);
FA fa2327(ip_55_16,ip_56_15,ip_57_14,p5830,p5831);
FA fa2328(ip_58_13,ip_59_12,ip_60_11,p5832,p5833);
FA fa2329(ip_61_10,ip_62_9,ip_63_8,p5834,p5835);
FA fa2330(p5642,p5644,p5660,p5836,p5837);
FA fa2331(p5670,p5672,p5678,p5838,p5839);
HA ha588(p5827,p5686,p5840,p5841);
FA fa2332(p5799,p5801,p5803,p5842,p5843);
FA fa2333(p5805,p5807,p5809,p5844,p5845);
FA fa2334(p5811,p5813,p5815,p5846,p5847);
FA fa2335(p5817,p5819,p5821,p5848,p5849);
FA fa2336(p5823,p5825,p5829,p5850,p5851);
FA fa2337(p5831,p5833,p5835,p5852,p5853);
FA fa2338(p5646,p5648,p5650,p5854,p5855);
FA fa2339(p5652,p5654,p5656,p5856,p5857);
FA fa2340(p5658,p5662,p5664,p5858,p5859);
FA fa2341(p5666,p5668,p5674,p5860,p5861);
HA ha589(p5676,p5680,p5862,p5863);
FA fa2342(p5682,p5696,p5698,p5864,p5865);
FA fa2343(p5702,p5704,p5837,p5866,p5867);
HA ha590(p5839,p5841,p5868,p5869);
FA fa2344(p5684,p5688,p5690,p5870,p5871);
FA fa2345(p5708,p5716,p5718,p5872,p5873);
FA fa2346(p5720,p5722,p5843,p5874,p5875);
FA fa2347(p5845,p5847,p5849,p5876,p5877);
HA ha591(p5851,p5853,p5878,p5879);
FA fa2348(p5863,p5869,p5692,p5880,p5881);
FA fa2349(p5694,p5700,p5728,p5882,p5883);
FA fa2350(p5855,p5857,p5859,p5884,p5885);
FA fa2351(p5861,p5865,p5867,p5886,p5887);
FA fa2352(p5879,p5706,p5710,p5888,p5889);
HA ha592(p5712,p5714,p5890,p5891);
FA fa2353(p5724,p5734,p5736,p5892,p5893);
FA fa2354(p5871,p5873,p5875,p5894,p5895);
FA fa2355(p5877,p5881,p5726,p5896,p5897);
FA fa2356(p5730,p5732,p5748,p5898,p5899);
HA ha593(p5750,p5883,p5900,p5901);
HA ha594(p5885,p5887,p5902,p5903);
FA fa2357(p5891,p5738,p5740,p5904,p5905);
FA fa2358(p5742,p5889,p5893,p5906,p5907);
FA fa2359(p5895,p5897,p5901,p5908,p5909);
FA fa2360(p5903,p5744,p5746,p5910,p5911);
HA ha595(p5752,p5899,p5912,p5913);
FA fa2361(p5754,p5756,p5905,p5914,p5915);
FA fa2362(p5907,p5909,p5913,p5916,p5917);
FA fa2363(p5758,p5760,p5762,p5918,p5919);
FA fa2364(p5772,p5911,p5764,p5920,p5921);
FA fa2365(p5766,p5915,p5917,p5922,p5923);
FA fa2366(p5768,p5770,p5919,p5924,p5925);
HA ha596(p5921,p5774,p5926,p5927);
FA fa2367(p5776,p5780,p5923,p5928,p5929);
FA fa2368(p5778,p5925,p5927,p5930,p5931);
HA ha597(p5929,p5782,p5932,p5933);
FA fa2369(p5784,p5931,p5933,p5934,p5935);
FA fa2370(p5786,p5788,p5935,p5936,p5937);
FA fa2371(p5790,p5937,p5794,p5938,p5939);
FA fa2372(p5792,p5939,p5796,p5940,p5941);
HA ha598(ip_9_63,ip_10_62,p5942,p5943);
FA fa2373(ip_11_61,ip_12_60,ip_13_59,p5944,p5945);
FA fa2374(ip_14_58,ip_15_57,ip_16_56,p5946,p5947);
FA fa2375(ip_17_55,ip_18_54,ip_19_53,p5948,p5949);
FA fa2376(ip_20_52,ip_21_51,ip_22_50,p5950,p5951);
HA ha599(ip_23_49,ip_24_48,p5952,p5953);
FA fa2377(ip_25_47,ip_26_46,ip_27_45,p5954,p5955);
FA fa2378(ip_28_44,ip_29_43,ip_30_42,p5956,p5957);
HA ha600(ip_31_41,ip_32_40,p5958,p5959);
HA ha601(ip_33_39,ip_34_38,p5960,p5961);
FA fa2379(ip_35_37,ip_36_36,ip_37_35,p5962,p5963);
FA fa2380(ip_38_34,ip_39_33,ip_40_32,p5964,p5965);
HA ha602(ip_41_31,ip_42_30,p5966,p5967);
FA fa2381(ip_43_29,ip_44_28,ip_45_27,p5968,p5969);
FA fa2382(ip_46_26,ip_47_25,ip_48_24,p5970,p5971);
FA fa2383(ip_49_23,ip_50_22,ip_51_21,p5972,p5973);
HA ha603(ip_52_20,ip_53_19,p5974,p5975);
FA fa2384(ip_54_18,ip_55_17,ip_56_16,p5976,p5977);
FA fa2385(ip_57_15,ip_58_14,ip_59_13,p5978,p5979);
FA fa2386(ip_60_12,ip_61_11,ip_62_10,p5980,p5981);
FA fa2387(ip_63_9,p5826,p5943,p5982,p5983);
FA fa2388(p5953,p5959,p5961,p5984,p5985);
FA fa2389(p5967,p5975,p5945,p5986,p5987);
FA fa2390(p5947,p5949,p5951,p5988,p5989);
FA fa2391(p5955,p5957,p5963,p5990,p5991);
HA ha604(p5965,p5969,p5992,p5993);
FA fa2392(p5971,p5973,p5977,p5994,p5995);
FA fa2393(p5979,p5981,p5798,p5996,p5997);
FA fa2394(p5800,p5802,p5804,p5998,p5999);
FA fa2395(p5806,p5808,p5810,p6000,p6001);
FA fa2396(p5812,p5814,p5816,p6002,p6003);
HA ha605(p5818,p5820,p6004,p6005);
FA fa2397(p5822,p5824,p5828,p6006,p6007);
FA fa2398(p5830,p5832,p5834,p6008,p6009);
FA fa2399(p5840,p5983,p5985,p6010,p6011);
FA fa2400(p5987,p5993,p5836,p6012,p6013);
FA fa2401(p5838,p5862,p5868,p6014,p6015);
FA fa2402(p5989,p5991,p5995,p6016,p6017);
FA fa2403(p5997,p6005,p5842,p6018,p6019);
FA fa2404(p5844,p5846,p5848,p6020,p6021);
FA fa2405(p5850,p5852,p5878,p6022,p6023);
FA fa2406(p5999,p6001,p6003,p6024,p6025);
FA fa2407(p6007,p6009,p6011,p6026,p6027);
FA fa2408(p6013,p5854,p5856,p6028,p6029);
FA fa2409(p5858,p5860,p5864,p6030,p6031);
FA fa2410(p5866,p6015,p6017,p6032,p6033);
FA fa2411(p6019,p5870,p5872,p6034,p6035);
FA fa2412(p5874,p5876,p5880,p6036,p6037);
HA ha606(p5890,p6021,p6038,p6039);
FA fa2413(p6023,p6025,p6027,p6040,p6041);
FA fa2414(p5882,p5884,p5886,p6042,p6043);
FA fa2415(p5900,p5902,p6029,p6044,p6045);
FA fa2416(p6031,p6033,p6039,p6046,p6047);
FA fa2417(p5888,p5892,p5894,p6048,p6049);
FA fa2418(p5896,p6035,p6037,p6050,p6051);
FA fa2419(p6041,p5898,p5912,p6052,p6053);
HA ha607(p6043,p6045,p6054,p6055);
FA fa2420(p6047,p5904,p5906,p6056,p6057);
FA fa2421(p5908,p6049,p6051,p6058,p6059);
FA fa2422(p6055,p5910,p6053,p6060,p6061);
FA fa2423(p5914,p5916,p6057,p6062,p6063);
FA fa2424(p6059,p5918,p5920,p6064,p6065);
FA fa2425(p6061,p5922,p5926,p6066,p6067);
FA fa2426(p6063,p5924,p6065,p6068,p6069);
FA fa2427(p5928,p6067,p5930,p6070,p6071);
FA fa2428(p5932,p6069,p6071,p6072,p6073);
FA fa2429(p5934,p6073,p5936,p6074,p6075);
FA fa2430(p6075,p5938,p5940,p6076,p6077);
FA fa2431(ip_10_63,ip_11_62,ip_12_61,p6078,p6079);
FA fa2432(ip_13_60,ip_14_59,ip_15_58,p6080,p6081);
FA fa2433(ip_16_57,ip_17_56,ip_18_55,p6082,p6083);
FA fa2434(ip_19_54,ip_20_53,ip_21_52,p6084,p6085);
FA fa2435(ip_22_51,ip_23_50,ip_24_49,p6086,p6087);
FA fa2436(ip_25_48,ip_26_47,ip_27_46,p6088,p6089);
FA fa2437(ip_28_45,ip_29_44,ip_30_43,p6090,p6091);
HA ha608(ip_31_42,ip_32_41,p6092,p6093);
FA fa2438(ip_33_40,ip_34_39,ip_35_38,p6094,p6095);
FA fa2439(ip_36_37,ip_37_36,ip_38_35,p6096,p6097);
FA fa2440(ip_39_34,ip_40_33,ip_41_32,p6098,p6099);
FA fa2441(ip_42_31,ip_43_30,ip_44_29,p6100,p6101);
HA ha609(ip_45_28,ip_46_27,p6102,p6103);
FA fa2442(ip_47_26,ip_48_25,ip_49_24,p6104,p6105);
HA ha610(ip_50_23,ip_51_22,p6106,p6107);
FA fa2443(ip_52_21,ip_53_20,ip_54_19,p6108,p6109);
FA fa2444(ip_55_18,ip_56_17,ip_57_16,p6110,p6111);
HA ha611(ip_58_15,ip_59_14,p6112,p6113);
FA fa2445(ip_60_13,ip_61_12,ip_62_11,p6114,p6115);
FA fa2446(ip_63_10,p5942,p5952,p6116,p6117);
HA ha612(p5958,p5960,p6118,p6119);
HA ha613(p5966,p5974,p6120,p6121);
FA fa2447(p6093,p6103,p6107,p6122,p6123);
FA fa2448(p6113,p6079,p6081,p6124,p6125);
HA ha614(p6083,p6085,p6126,p6127);
HA ha615(p6087,p6089,p6128,p6129);
HA ha616(p6091,p6095,p6130,p6131);
HA ha617(p6097,p6099,p6132,p6133);
FA fa2449(p6101,p6105,p6109,p6134,p6135);
FA fa2450(p6111,p6115,p6119,p6136,p6137);
FA fa2451(p6121,p5944,p5946,p6138,p6139);
HA ha618(p5948,p5950,p6140,p6141);
FA fa2452(p5954,p5956,p5962,p6142,p6143);
HA ha619(p5964,p5968,p6144,p6145);
FA fa2453(p5970,p5972,p5976,p6146,p6147);
FA fa2454(p5978,p5980,p5992,p6148,p6149);
HA ha620(p6117,p6123,p6150,p6151);
HA ha621(p6127,p6129,p6152,p6153);
HA ha622(p6131,p6133,p6154,p6155);
FA fa2455(p5982,p5984,p5986,p6156,p6157);
FA fa2456(p6004,p6125,p6135,p6158,p6159);
FA fa2457(p6137,p6141,p6145,p6160,p6161);
FA fa2458(p6151,p6153,p6155,p6162,p6163);
HA ha623(p5988,p5990,p6164,p6165);
FA fa2459(p5994,p5996,p6139,p6166,p6167);
FA fa2460(p6143,p6147,p6149,p6168,p6169);
FA fa2461(p5998,p6000,p6002,p6170,p6171);
HA ha624(p6006,p6008,p6172,p6173);
FA fa2462(p6010,p6012,p6157,p6174,p6175);
FA fa2463(p6159,p6161,p6163,p6176,p6177);
FA fa2464(p6165,p6014,p6016,p6178,p6179);
FA fa2465(p6018,p6167,p6169,p6180,p6181);
FA fa2466(p6173,p6020,p6022,p6182,p6183);
FA fa2467(p6024,p6026,p6038,p6184,p6185);
FA fa2468(p6171,p6175,p6177,p6186,p6187);
FA fa2469(p6028,p6030,p6032,p6188,p6189);
HA ha625(p6179,p6181,p6190,p6191);
FA fa2470(p6034,p6036,p6040,p6192,p6193);
FA fa2471(p6183,p6185,p6187,p6194,p6195);
FA fa2472(p6191,p6042,p6044,p6196,p6197);
FA fa2473(p6046,p6054,p6189,p6198,p6199);
FA fa2474(p6048,p6050,p6193,p6200,p6201);
FA fa2475(p6195,p6052,p6197,p6202,p6203);
FA fa2476(p6199,p6056,p6058,p6204,p6205);
FA fa2477(p6201,p6060,p6203,p6206,p6207);
FA fa2478(p6062,p6205,p6064,p6208,p6209);
FA fa2479(p6207,p6066,p6209,p6210,p6211);
FA fa2480(p6068,p6070,p6211,p6212,p6213);
FA fa2481(p6072,p6213,p6074,p6214,p6215);
HA ha626(ip_11_63,ip_12_62,p6216,p6217);
FA fa2482(ip_13_61,ip_14_60,ip_15_59,p6218,p6219);
FA fa2483(ip_16_58,ip_17_57,ip_18_56,p6220,p6221);
FA fa2484(ip_19_55,ip_20_54,ip_21_53,p6222,p6223);
FA fa2485(ip_22_52,ip_23_51,ip_24_50,p6224,p6225);
FA fa2486(ip_25_49,ip_26_48,ip_27_47,p6226,p6227);
FA fa2487(ip_28_46,ip_29_45,ip_30_44,p6228,p6229);
FA fa2488(ip_31_43,ip_32_42,ip_33_41,p6230,p6231);
FA fa2489(ip_34_40,ip_35_39,ip_36_38,p6232,p6233);
FA fa2490(ip_37_37,ip_38_36,ip_39_35,p6234,p6235);
FA fa2491(ip_40_34,ip_41_33,ip_42_32,p6236,p6237);
FA fa2492(ip_43_31,ip_44_30,ip_45_29,p6238,p6239);
FA fa2493(ip_46_28,ip_47_27,ip_48_26,p6240,p6241);
FA fa2494(ip_49_25,ip_50_24,ip_51_23,p6242,p6243);
HA ha627(ip_52_22,ip_53_21,p6244,p6245);
HA ha628(ip_54_20,ip_55_19,p6246,p6247);
FA fa2495(ip_56_18,ip_57_17,ip_58_16,p6248,p6249);
FA fa2496(ip_59_15,ip_60_14,ip_61_13,p6250,p6251);
FA fa2497(ip_62_12,ip_63_11,p6092,p6252,p6253);
FA fa2498(p6102,p6106,p6112,p6254,p6255);
FA fa2499(p6217,p6245,p6247,p6256,p6257);
FA fa2500(p6118,p6120,p6219,p6258,p6259);
FA fa2501(p6221,p6223,p6225,p6260,p6261);
FA fa2502(p6227,p6229,p6231,p6262,p6263);
FA fa2503(p6233,p6235,p6237,p6264,p6265);
FA fa2504(p6239,p6241,p6243,p6266,p6267);
FA fa2505(p6249,p6251,p6253,p6268,p6269);
HA ha629(p6078,p6080,p6270,p6271);
HA ha630(p6082,p6084,p6272,p6273);
FA fa2506(p6086,p6088,p6090,p6274,p6275);
HA ha631(p6094,p6096,p6276,p6277);
FA fa2507(p6098,p6100,p6104,p6278,p6279);
FA fa2508(p6108,p6110,p6114,p6280,p6281);
FA fa2509(p6126,p6128,p6130,p6282,p6283);
HA ha632(p6132,p6255,p6284,p6285);
FA fa2510(p6257,p6116,p6122,p6286,p6287);
FA fa2511(p6140,p6144,p6150,p6288,p6289);
FA fa2512(p6152,p6154,p6259,p6290,p6291);
FA fa2513(p6261,p6263,p6265,p6292,p6293);
FA fa2514(p6267,p6269,p6271,p6294,p6295);
FA fa2515(p6273,p6277,p6285,p6296,p6297);
HA ha633(p6124,p6134,p6298,p6299);
FA fa2516(p6136,p6275,p6279,p6300,p6301);
FA fa2517(p6281,p6283,p6138,p6302,p6303);
FA fa2518(p6142,p6146,p6148,p6304,p6305);
HA ha634(p6164,p6287,p6306,p6307);
HA ha635(p6289,p6291,p6308,p6309);
HA ha636(p6293,p6295,p6310,p6311);
FA fa2519(p6297,p6299,p6156,p6312,p6313);
HA ha637(p6158,p6160,p6314,p6315);
HA ha638(p6162,p6172,p6316,p6317);
HA ha639(p6301,p6303,p6318,p6319);
FA fa2520(p6307,p6309,p6311,p6320,p6321);
FA fa2521(p6166,p6168,p6305,p6322,p6323);
FA fa2522(p6313,p6315,p6317,p6324,p6325);
FA fa2523(p6319,p6170,p6174,p6326,p6327);
FA fa2524(p6176,p6321,p6178,p6328,p6329);
FA fa2525(p6180,p6190,p6323,p6330,p6331);
FA fa2526(p6325,p6182,p6184,p6332,p6333);
FA fa2527(p6186,p6327,p6329,p6334,p6335);
FA fa2528(p6188,p6331,p6192,p6336,p6337);
FA fa2529(p6194,p6333,p6335,p6338,p6339);
FA fa2530(p6196,p6198,p6337,p6340,p6341);
FA fa2531(p6200,p6339,p6202,p6342,p6343);
FA fa2532(p6341,p6204,p6343,p6344,p6345);
FA fa2533(p6206,p6208,p6345,p6346,p6347);
FA fa2534(p6210,p6347,p6212,p6348,p6349);
FA fa2535(ip_12_63,ip_13_62,ip_14_61,p6350,p6351);
HA ha640(ip_15_60,ip_16_59,p6352,p6353);
FA fa2536(ip_17_58,ip_18_57,ip_19_56,p6354,p6355);
FA fa2537(ip_20_55,ip_21_54,ip_22_53,p6356,p6357);
FA fa2538(ip_23_52,ip_24_51,ip_25_50,p6358,p6359);
HA ha641(ip_26_49,ip_27_48,p6360,p6361);
FA fa2539(ip_28_47,ip_29_46,ip_30_45,p6362,p6363);
FA fa2540(ip_31_44,ip_32_43,ip_33_42,p6364,p6365);
FA fa2541(ip_34_41,ip_35_40,ip_36_39,p6366,p6367);
FA fa2542(ip_37_38,ip_38_37,ip_39_36,p6368,p6369);
FA fa2543(ip_40_35,ip_41_34,ip_42_33,p6370,p6371);
HA ha642(ip_43_32,ip_44_31,p6372,p6373);
FA fa2544(ip_45_30,ip_46_29,ip_47_28,p6374,p6375);
FA fa2545(ip_48_27,ip_49_26,ip_50_25,p6376,p6377);
FA fa2546(ip_51_24,ip_52_23,ip_53_22,p6378,p6379);
FA fa2547(ip_54_21,ip_55_20,ip_56_19,p6380,p6381);
FA fa2548(ip_57_18,ip_58_17,ip_59_16,p6382,p6383);
FA fa2549(ip_60_15,ip_61_14,ip_62_13,p6384,p6385);
FA fa2550(ip_63_12,p6216,p6244,p6386,p6387);
FA fa2551(p6246,p6353,p6361,p6388,p6389);
FA fa2552(p6373,p6351,p6355,p6390,p6391);
FA fa2553(p6357,p6359,p6363,p6392,p6393);
HA ha643(p6365,p6367,p6394,p6395);
FA fa2554(p6369,p6371,p6375,p6396,p6397);
FA fa2555(p6377,p6379,p6381,p6398,p6399);
FA fa2556(p6383,p6385,p6218,p6400,p6401);
FA fa2557(p6220,p6222,p6224,p6402,p6403);
FA fa2558(p6226,p6228,p6230,p6404,p6405);
FA fa2559(p6232,p6234,p6236,p6406,p6407);
FA fa2560(p6238,p6240,p6242,p6408,p6409);
FA fa2561(p6248,p6250,p6252,p6410,p6411);
FA fa2562(p6387,p6389,p6395,p6412,p6413);
FA fa2563(p6254,p6256,p6270,p6414,p6415);
FA fa2564(p6272,p6276,p6284,p6416,p6417);
FA fa2565(p6391,p6393,p6397,p6418,p6419);
FA fa2566(p6399,p6401,p6258,p6420,p6421);
FA fa2567(p6260,p6262,p6264,p6422,p6423);
HA ha644(p6266,p6268,p6424,p6425);
FA fa2568(p6403,p6405,p6407,p6426,p6427);
HA ha645(p6409,p6411,p6428,p6429);
FA fa2569(p6413,p6274,p6278,p6430,p6431);
HA ha646(p6280,p6282,p6432,p6433);
FA fa2570(p6298,p6415,p6417,p6434,p6435);
HA ha647(p6419,p6421,p6436,p6437);
FA fa2571(p6425,p6429,p6286,p6438,p6439);
FA fa2572(p6288,p6290,p6292,p6440,p6441);
FA fa2573(p6294,p6296,p6306,p6442,p6443);
FA fa2574(p6308,p6310,p6423,p6444,p6445);
HA ha648(p6427,p6433,p6446,p6447);
FA fa2575(p6437,p6300,p6302,p6448,p6449);
FA fa2576(p6314,p6316,p6318,p6450,p6451);
FA fa2577(p6431,p6435,p6439,p6452,p6453);
FA fa2578(p6447,p6304,p6312,p6454,p6455);
HA ha649(p6441,p6443,p6456,p6457);
FA fa2579(p6445,p6320,p6449,p6458,p6459);
HA ha650(p6451,p6453,p6460,p6461);
FA fa2580(p6457,p6322,p6324,p6462,p6463);
FA fa2581(p6455,p6461,p6326,p6464,p6465);
FA fa2582(p6328,p6459,p6330,p6466,p6467);
FA fa2583(p6463,p6465,p6332,p6468,p6469);
HA ha651(p6334,p6467,p6470,p6471);
FA fa2584(p6336,p6469,p6471,p6472,p6473);
FA fa2585(p6338,p6340,p6473,p6474,p6475);
FA fa2586(p6342,p6475,p6344,p6476,p6477);
FA fa2587(p6477,p6346,p6348,p6478,p6479);
FA fa2588(ip_13_63,ip_14_62,ip_15_61,p6480,p6481);
FA fa2589(ip_16_60,ip_17_59,ip_18_58,p6482,p6483);
FA fa2590(ip_19_57,ip_20_56,ip_21_55,p6484,p6485);
FA fa2591(ip_22_54,ip_23_53,ip_24_52,p6486,p6487);
HA ha652(ip_25_51,ip_26_50,p6488,p6489);
FA fa2592(ip_27_49,ip_28_48,ip_29_47,p6490,p6491);
FA fa2593(ip_30_46,ip_31_45,ip_32_44,p6492,p6493);
HA ha653(ip_33_43,ip_34_42,p6494,p6495);
FA fa2594(ip_35_41,ip_36_40,ip_37_39,p6496,p6497);
FA fa2595(ip_38_38,ip_39_37,ip_40_36,p6498,p6499);
HA ha654(ip_41_35,ip_42_34,p6500,p6501);
HA ha655(ip_43_33,ip_44_32,p6502,p6503);
HA ha656(ip_45_31,ip_46_30,p6504,p6505);
FA fa2596(ip_47_29,ip_48_28,ip_49_27,p6506,p6507);
HA ha657(ip_50_26,ip_51_25,p6508,p6509);
HA ha658(ip_52_24,ip_53_23,p6510,p6511);
FA fa2597(ip_54_22,ip_55_21,ip_56_20,p6512,p6513);
FA fa2598(ip_57_19,ip_58_18,ip_59_17,p6514,p6515);
FA fa2599(ip_60_16,ip_61_15,ip_62_14,p6516,p6517);
FA fa2600(ip_63_13,p6352,p6360,p6518,p6519);
FA fa2601(p6372,p6489,p6495,p6520,p6521);
FA fa2602(p6501,p6503,p6505,p6522,p6523);
FA fa2603(p6509,p6511,p6481,p6524,p6525);
FA fa2604(p6483,p6485,p6487,p6526,p6527);
FA fa2605(p6491,p6493,p6497,p6528,p6529);
HA ha659(p6499,p6507,p6530,p6531);
FA fa2606(p6513,p6515,p6517,p6532,p6533);
FA fa2607(p6350,p6354,p6356,p6534,p6535);
FA fa2608(p6358,p6362,p6364,p6536,p6537);
FA fa2609(p6366,p6368,p6370,p6538,p6539);
FA fa2610(p6374,p6376,p6378,p6540,p6541);
HA ha660(p6380,p6382,p6542,p6543);
HA ha661(p6384,p6394,p6544,p6545);
HA ha662(p6519,p6521,p6546,p6547);
FA fa2611(p6523,p6525,p6531,p6548,p6549);
HA ha663(p6386,p6388,p6550,p6551);
FA fa2612(p6527,p6529,p6533,p6552,p6553);
FA fa2613(p6543,p6545,p6547,p6554,p6555);
FA fa2614(p6390,p6392,p6396,p6556,p6557);
HA ha664(p6398,p6400,p6558,p6559);
FA fa2615(p6535,p6537,p6539,p6560,p6561);
FA fa2616(p6541,p6549,p6551,p6562,p6563);
FA fa2617(p6402,p6404,p6406,p6564,p6565);
HA ha665(p6408,p6410,p6566,p6567);
FA fa2618(p6412,p6424,p6428,p6568,p6569);
FA fa2619(p6553,p6555,p6559,p6570,p6571);
HA ha666(p6414,p6416,p6572,p6573);
HA ha667(p6418,p6420,p6574,p6575);
HA ha668(p6432,p6436,p6576,p6577);
FA fa2620(p6557,p6561,p6563,p6578,p6579);
FA fa2621(p6567,p6422,p6426,p6580,p6581);
FA fa2622(p6446,p6565,p6569,p6582,p6583);
FA fa2623(p6571,p6573,p6575,p6584,p6585);
FA fa2624(p6577,p6430,p6434,p6586,p6587);
FA fa2625(p6438,p6579,p6440,p6588,p6589);
FA fa2626(p6442,p6444,p6456,p6590,p6591);
FA fa2627(p6581,p6583,p6585,p6592,p6593);
HA ha669(p6448,p6450,p6594,p6595);
FA fa2628(p6452,p6460,p6587,p6596,p6597);
FA fa2629(p6589,p6454,p6591,p6598,p6599);
FA fa2630(p6593,p6595,p6458,p6600,p6601);
FA fa2631(p6597,p6462,p6464,p6602,p6603);
FA fa2632(p6599,p6601,p6466,p6604,p6605);
FA fa2633(p6470,p6468,p6603,p6606,p6607);
FA fa2634(p6605,p6472,p6607,p6608,p6609);
FA fa2635(p6474,p6609,p6476,p6610,p6611);
FA fa2636(ip_14_63,ip_15_62,ip_16_61,p6612,p6613);
FA fa2637(ip_17_60,ip_18_59,ip_19_58,p6614,p6615);
FA fa2638(ip_20_57,ip_21_56,ip_22_55,p6616,p6617);
HA ha670(ip_23_54,ip_24_53,p6618,p6619);
FA fa2639(ip_25_52,ip_26_51,ip_27_50,p6620,p6621);
HA ha671(ip_28_49,ip_29_48,p6622,p6623);
HA ha672(ip_30_47,ip_31_46,p6624,p6625);
FA fa2640(ip_32_45,ip_33_44,ip_34_43,p6626,p6627);
FA fa2641(ip_35_42,ip_36_41,ip_37_40,p6628,p6629);
FA fa2642(ip_38_39,ip_39_38,ip_40_37,p6630,p6631);
FA fa2643(ip_41_36,ip_42_35,ip_43_34,p6632,p6633);
HA ha673(ip_44_33,ip_45_32,p6634,p6635);
FA fa2644(ip_46_31,ip_47_30,ip_48_29,p6636,p6637);
FA fa2645(ip_49_28,ip_50_27,ip_51_26,p6638,p6639);
HA ha674(ip_52_25,ip_53_24,p6640,p6641);
FA fa2646(ip_54_23,ip_55_22,ip_56_21,p6642,p6643);
FA fa2647(ip_57_20,ip_58_19,ip_59_18,p6644,p6645);
FA fa2648(ip_60_17,ip_61_16,ip_62_15,p6646,p6647);
FA fa2649(ip_63_14,p6488,p6494,p6648,p6649);
FA fa2650(p6500,p6502,p6504,p6650,p6651);
FA fa2651(p6508,p6510,p6619,p6652,p6653);
FA fa2652(p6623,p6625,p6635,p6654,p6655);
HA ha675(p6641,p6613,p6656,p6657);
FA fa2653(p6615,p6617,p6621,p6658,p6659);
FA fa2654(p6627,p6629,p6631,p6660,p6661);
HA ha676(p6633,p6637,p6662,p6663);
FA fa2655(p6639,p6643,p6645,p6664,p6665);
HA ha677(p6647,p6480,p6666,p6667);
FA fa2656(p6482,p6484,p6486,p6668,p6669);
FA fa2657(p6490,p6492,p6496,p6670,p6671);
FA fa2658(p6498,p6506,p6512,p6672,p6673);
FA fa2659(p6514,p6516,p6530,p6674,p6675);
FA fa2660(p6649,p6651,p6653,p6676,p6677);
HA ha678(p6655,p6657,p6678,p6679);
FA fa2661(p6663,p6518,p6520,p6680,p6681);
FA fa2662(p6522,p6524,p6542,p6682,p6683);
FA fa2663(p6544,p6546,p6659,p6684,p6685);
FA fa2664(p6661,p6665,p6667,p6686,p6687);
FA fa2665(p6679,p6526,p6528,p6688,p6689);
FA fa2666(p6532,p6550,p6669,p6690,p6691);
FA fa2667(p6671,p6673,p6675,p6692,p6693);
FA fa2668(p6677,p6534,p6536,p6694,p6695);
FA fa2669(p6538,p6540,p6548,p6696,p6697);
FA fa2670(p6558,p6681,p6683,p6698,p6699);
FA fa2671(p6685,p6687,p6552,p6700,p6701);
FA fa2672(p6554,p6566,p6689,p6702,p6703);
FA fa2673(p6691,p6693,p6556,p6704,p6705);
FA fa2674(p6560,p6562,p6572,p6706,p6707);
HA ha679(p6574,p6576,p6708,p6709);
FA fa2675(p6695,p6697,p6699,p6710,p6711);
FA fa2676(p6701,p6564,p6568,p6712,p6713);
FA fa2677(p6570,p6703,p6705,p6714,p6715);
HA ha680(p6709,p6578,p6716,p6717);
FA fa2678(p6707,p6711,p6580,p6718,p6719);
FA fa2679(p6582,p6584,p6713,p6720,p6721);
FA fa2680(p6715,p6717,p6586,p6722,p6723);
FA fa2681(p6588,p6594,p6719,p6724,p6725);
FA fa2682(p6590,p6592,p6721,p6726,p6727);
FA fa2683(p6723,p6596,p6725,p6728,p6729);
FA fa2684(p6598,p6600,p6727,p6730,p6731);
FA fa2685(p6729,p6602,p6604,p6732,p6733);
FA fa2686(p6731,p6606,p6733,p6734,p6735);
FA fa2687(p6608,p6735,p6610,p6736,p6737);
FA fa2688(ip_15_63,ip_16_62,ip_17_61,p6738,p6739);
HA ha681(ip_18_60,ip_19_59,p6740,p6741);
FA fa2689(ip_20_58,ip_21_57,ip_22_56,p6742,p6743);
FA fa2690(ip_23_55,ip_24_54,ip_25_53,p6744,p6745);
FA fa2691(ip_26_52,ip_27_51,ip_28_50,p6746,p6747);
FA fa2692(ip_29_49,ip_30_48,ip_31_47,p6748,p6749);
FA fa2693(ip_32_46,ip_33_45,ip_34_44,p6750,p6751);
FA fa2694(ip_35_43,ip_36_42,ip_37_41,p6752,p6753);
FA fa2695(ip_38_40,ip_39_39,ip_40_38,p6754,p6755);
FA fa2696(ip_41_37,ip_42_36,ip_43_35,p6756,p6757);
FA fa2697(ip_44_34,ip_45_33,ip_46_32,p6758,p6759);
FA fa2698(ip_47_31,ip_48_30,ip_49_29,p6760,p6761);
HA ha682(ip_50_28,ip_51_27,p6762,p6763);
FA fa2699(ip_52_26,ip_53_25,ip_54_24,p6764,p6765);
FA fa2700(ip_55_23,ip_56_22,ip_57_21,p6766,p6767);
HA ha683(ip_58_20,ip_59_19,p6768,p6769);
FA fa2701(ip_60_18,ip_61_17,ip_62_16,p6770,p6771);
FA fa2702(ip_63_15,p6618,p6622,p6772,p6773);
FA fa2703(p6624,p6634,p6640,p6774,p6775);
FA fa2704(p6741,p6763,p6769,p6776,p6777);
FA fa2705(p6739,p6743,p6745,p6778,p6779);
FA fa2706(p6747,p6749,p6751,p6780,p6781);
FA fa2707(p6753,p6755,p6757,p6782,p6783);
HA ha684(p6759,p6761,p6784,p6785);
FA fa2708(p6765,p6767,p6771,p6786,p6787);
HA ha685(p6612,p6614,p6788,p6789);
HA ha686(p6616,p6620,p6790,p6791);
FA fa2709(p6626,p6628,p6630,p6792,p6793);
FA fa2710(p6632,p6636,p6638,p6794,p6795);
HA ha687(p6642,p6644,p6796,p6797);
FA fa2711(p6646,p6656,p6662,p6798,p6799);
FA fa2712(p6773,p6775,p6777,p6800,p6801);
FA fa2713(p6785,p6648,p6650,p6802,p6803);
HA ha688(p6652,p6654,p6804,p6805);
FA fa2714(p6666,p6678,p6779,p6806,p6807);
HA ha689(p6781,p6783,p6808,p6809);
FA fa2715(p6787,p6789,p6791,p6810,p6811);
FA fa2716(p6797,p6658,p6660,p6812,p6813);
FA fa2717(p6664,p6793,p6795,p6814,p6815);
FA fa2718(p6799,p6801,p6805,p6816,p6817);
FA fa2719(p6809,p6668,p6670,p6818,p6819);
FA fa2720(p6672,p6674,p6676,p6820,p6821);
FA fa2721(p6803,p6807,p6811,p6822,p6823);
FA fa2722(p6680,p6682,p6684,p6824,p6825);
HA ha690(p6686,p6813,p6826,p6827);
HA ha691(p6815,p6817,p6828,p6829);
FA fa2723(p6688,p6690,p6692,p6830,p6831);
FA fa2724(p6819,p6821,p6823,p6832,p6833);
HA ha692(p6827,p6829,p6834,p6835);
HA ha693(p6694,p6696,p6836,p6837);
FA fa2725(p6698,p6700,p6708,p6838,p6839);
HA ha694(p6825,p6835,p6840,p6841);
HA ha695(p6702,p6704,p6842,p6843);
HA ha696(p6831,p6833,p6844,p6845);
FA fa2726(p6837,p6841,p6706,p6846,p6847);
FA fa2727(p6710,p6716,p6839,p6848,p6849);
FA fa2728(p6843,p6845,p6712,p6850,p6851);
FA fa2729(p6714,p6847,p6718,p6852,p6853);
FA fa2730(p6849,p6851,p6720,p6854,p6855);
HA ha697(p6722,p6853,p6856,p6857);
HA ha698(p6724,p6855,p6858,p6859);
FA fa2731(p6857,p6726,p6859,p6860,p6861);
FA fa2732(p6728,p6730,p6861,p6862,p6863);
HA ha699(p6732,p6863,p6864,p6865);
HA ha700(p6865,p6734,p6866,p6867);
HA ha701(ip_16_63,ip_17_62,p6868,p6869);
FA fa2733(ip_18_61,ip_19_60,ip_20_59,p6870,p6871);
FA fa2734(ip_21_58,ip_22_57,ip_23_56,p6872,p6873);
FA fa2735(ip_24_55,ip_25_54,ip_26_53,p6874,p6875);
FA fa2736(ip_27_52,ip_28_51,ip_29_50,p6876,p6877);
FA fa2737(ip_30_49,ip_31_48,ip_32_47,p6878,p6879);
FA fa2738(ip_33_46,ip_34_45,ip_35_44,p6880,p6881);
FA fa2739(ip_36_43,ip_37_42,ip_38_41,p6882,p6883);
FA fa2740(ip_39_40,ip_40_39,ip_41_38,p6884,p6885);
FA fa2741(ip_42_37,ip_43_36,ip_44_35,p6886,p6887);
FA fa2742(ip_45_34,ip_46_33,ip_47_32,p6888,p6889);
FA fa2743(ip_48_31,ip_49_30,ip_50_29,p6890,p6891);
HA ha702(ip_51_28,ip_52_27,p6892,p6893);
FA fa2744(ip_53_26,ip_54_25,ip_55_24,p6894,p6895);
FA fa2745(ip_56_23,ip_57_22,ip_58_21,p6896,p6897);
FA fa2746(ip_59_20,ip_60_19,ip_61_18,p6898,p6899);
FA fa2747(ip_62_17,ip_63_16,p6740,p6900,p6901);
FA fa2748(p6762,p6768,p6869,p6902,p6903);
FA fa2749(p6893,p6871,p6873,p6904,p6905);
FA fa2750(p6875,p6877,p6879,p6906,p6907);
FA fa2751(p6881,p6883,p6885,p6908,p6909);
FA fa2752(p6887,p6889,p6891,p6910,p6911);
FA fa2753(p6895,p6897,p6899,p6912,p6913);
HA ha703(p6901,p6738,p6914,p6915);
FA fa2754(p6742,p6744,p6746,p6916,p6917);
HA ha704(p6748,p6750,p6918,p6919);
FA fa2755(p6752,p6754,p6756,p6920,p6921);
FA fa2756(p6758,p6760,p6764,p6922,p6923);
HA ha705(p6766,p6770,p6924,p6925);
FA fa2757(p6784,p6903,p6772,p6926,p6927);
FA fa2758(p6774,p6776,p6788,p6928,p6929);
FA fa2759(p6790,p6796,p6905,p6930,p6931);
HA ha706(p6907,p6909,p6932,p6933);
HA ha707(p6911,p6913,p6934,p6935);
FA fa2760(p6915,p6919,p6925,p6936,p6937);
FA fa2761(p6778,p6780,p6782,p6938,p6939);
FA fa2762(p6786,p6804,p6808,p6940,p6941);
FA fa2763(p6917,p6921,p6923,p6942,p6943);
FA fa2764(p6927,p6933,p6935,p6944,p6945);
FA fa2765(p6792,p6794,p6798,p6946,p6947);
FA fa2766(p6800,p6929,p6931,p6948,p6949);
FA fa2767(p6937,p6802,p6806,p6950,p6951);
FA fa2768(p6810,p6939,p6941,p6952,p6953);
HA ha708(p6943,p6945,p6954,p6955);
FA fa2769(p6812,p6814,p6816,p6956,p6957);
FA fa2770(p6826,p6828,p6947,p6958,p6959);
FA fa2771(p6949,p6955,p6818,p6960,p6961);
HA ha709(p6820,p6822,p6962,p6963);
FA fa2772(p6834,p6951,p6953,p6964,p6965);
FA fa2773(p6824,p6836,p6840,p6966,p6967);
FA fa2774(p6957,p6959,p6961,p6968,p6969);
FA fa2775(p6963,p6830,p6832,p6970,p6971);
HA ha710(p6842,p6844,p6972,p6973);
FA fa2776(p6965,p6838,p6967,p6974,p6975);
FA fa2777(p6969,p6973,p6846,p6976,p6977);
FA fa2778(p6971,p6848,p6850,p6978,p6979);
FA fa2779(p6975,p6977,p6852,p6980,p6981);
FA fa2780(p6856,p6854,p6858,p6982,p6983);
FA fa2781(p6979,p6981,p6983,p6984,p6985);
FA fa2782(p6860,p6985,p6862,p6986,p6987);
FA fa2783(p6864,p6987,p6866,p6988,p6989);
FA fa2784(ip_17_63,ip_18_62,ip_19_61,p6990,p6991);
FA fa2785(ip_20_60,ip_21_59,ip_22_58,p6992,p6993);
FA fa2786(ip_23_57,ip_24_56,ip_25_55,p6994,p6995);
FA fa2787(ip_26_54,ip_27_53,ip_28_52,p6996,p6997);
FA fa2788(ip_29_51,ip_30_50,ip_31_49,p6998,p6999);
HA ha711(ip_32_48,ip_33_47,p7000,p7001);
FA fa2789(ip_34_46,ip_35_45,ip_36_44,p7002,p7003);
HA ha712(ip_37_43,ip_38_42,p7004,p7005);
HA ha713(ip_39_41,ip_40_40,p7006,p7007);
FA fa2790(ip_41_39,ip_42_38,ip_43_37,p7008,p7009);
FA fa2791(ip_44_36,ip_45_35,ip_46_34,p7010,p7011);
HA ha714(ip_47_33,ip_48_32,p7012,p7013);
FA fa2792(ip_49_31,ip_50_30,ip_51_29,p7014,p7015);
FA fa2793(ip_52_28,ip_53_27,ip_54_26,p7016,p7017);
FA fa2794(ip_55_25,ip_56_24,ip_57_23,p7018,p7019);
FA fa2795(ip_58_22,ip_59_21,ip_60_20,p7020,p7021);
FA fa2796(ip_61_19,ip_62_18,ip_63_17,p7022,p7023);
FA fa2797(p6868,p6892,p7001,p7024,p7025);
HA ha715(p7005,p7007,p7026,p7027);
HA ha716(p7013,p6991,p7028,p7029);
FA fa2798(p6993,p6995,p6997,p7030,p7031);
FA fa2799(p6999,p7003,p7009,p7032,p7033);
FA fa2800(p7011,p7015,p7017,p7034,p7035);
FA fa2801(p7019,p7021,p7023,p7036,p7037);
FA fa2802(p7027,p6870,p6872,p7038,p7039);
FA fa2803(p6874,p6876,p6878,p7040,p7041);
FA fa2804(p6880,p6882,p6884,p7042,p7043);
FA fa2805(p6886,p6888,p6890,p7044,p7045);
FA fa2806(p6894,p6896,p6898,p7046,p7047);
HA ha717(p6900,p7025,p7048,p7049);
FA fa2807(p7029,p6902,p6914,p7050,p7051);
FA fa2808(p6918,p6924,p7031,p7052,p7053);
FA fa2809(p7033,p7035,p7037,p7054,p7055);
HA ha718(p7049,p6904,p7056,p7057);
FA fa2810(p6906,p6908,p6910,p7058,p7059);
FA fa2811(p6912,p6932,p6934,p7060,p7061);
FA fa2812(p7039,p7041,p7043,p7062,p7063);
HA ha719(p7045,p7047,p7064,p7065);
FA fa2813(p6916,p6920,p6922,p7066,p7067);
FA fa2814(p6926,p7051,p7053,p7068,p7069);
FA fa2815(p7055,p7057,p7065,p7070,p7071);
FA fa2816(p6928,p6930,p6936,p7072,p7073);
FA fa2817(p7059,p7061,p7063,p7074,p7075);
FA fa2818(p6938,p6940,p6942,p7076,p7077);
FA fa2819(p6944,p6954,p7067,p7078,p7079);
FA fa2820(p7069,p7071,p6946,p7080,p7081);
HA ha720(p6948,p7073,p7082,p7083);
FA fa2821(p7075,p6950,p6952,p7084,p7085);
FA fa2822(p6962,p7077,p7079,p7086,p7087);
FA fa2823(p7081,p7083,p6956,p7088,p7089);
FA fa2824(p6958,p6960,p6964,p7090,p7091);
FA fa2825(p6972,p7085,p7087,p7092,p7093);
HA ha721(p7089,p6966,p7094,p7095);
HA ha722(p6968,p7091,p7096,p7097);
FA fa2826(p6970,p7093,p7095,p7098,p7099);
FA fa2827(p7097,p6974,p6976,p7100,p7101);
FA fa2828(p7099,p6978,p6980,p7102,p7103);
FA fa2829(p7101,p6982,p7103,p7104,p7105);
FA fa2830(p6984,p7105,p6986,p7106,p7107);
FA fa2831(ip_18_63,ip_19_62,ip_20_61,p7108,p7109);
FA fa2832(ip_21_60,ip_22_59,ip_23_58,p7110,p7111);
FA fa2833(ip_24_57,ip_25_56,ip_26_55,p7112,p7113);
FA fa2834(ip_27_54,ip_28_53,ip_29_52,p7114,p7115);
FA fa2835(ip_30_51,ip_31_50,ip_32_49,p7116,p7117);
HA ha723(ip_33_48,ip_34_47,p7118,p7119);
FA fa2836(ip_35_46,ip_36_45,ip_37_44,p7120,p7121);
FA fa2837(ip_38_43,ip_39_42,ip_40_41,p7122,p7123);
HA ha724(ip_41_40,ip_42_39,p7124,p7125);
FA fa2838(ip_43_38,ip_44_37,ip_45_36,p7126,p7127);
FA fa2839(ip_46_35,ip_47_34,ip_48_33,p7128,p7129);
FA fa2840(ip_49_32,ip_50_31,ip_51_30,p7130,p7131);
FA fa2841(ip_52_29,ip_53_28,ip_54_27,p7132,p7133);
FA fa2842(ip_55_26,ip_56_25,ip_57_24,p7134,p7135);
FA fa2843(ip_58_23,ip_59_22,ip_60_21,p7136,p7137);
FA fa2844(ip_61_20,ip_62_19,ip_63_18,p7138,p7139);
FA fa2845(p7000,p7004,p7006,p7140,p7141);
HA ha725(p7012,p7119,p7142,p7143);
FA fa2846(p7125,p7026,p7109,p7144,p7145);
FA fa2847(p7111,p7113,p7115,p7146,p7147);
FA fa2848(p7117,p7121,p7123,p7148,p7149);
FA fa2849(p7127,p7129,p7131,p7150,p7151);
FA fa2850(p7133,p7135,p7137,p7152,p7153);
FA fa2851(p7139,p7143,p6990,p7154,p7155);
FA fa2852(p6992,p6994,p6996,p7156,p7157);
FA fa2853(p6998,p7002,p7008,p7158,p7159);
FA fa2854(p7010,p7014,p7016,p7160,p7161);
FA fa2855(p7018,p7020,p7022,p7162,p7163);
FA fa2856(p7028,p7141,p7024,p7164,p7165);
HA ha726(p7048,p7145,p7166,p7167);
FA fa2857(p7147,p7149,p7151,p7168,p7169);
FA fa2858(p7153,p7155,p7030,p7170,p7171);
FA fa2859(p7032,p7034,p7036,p7172,p7173);
FA fa2860(p7157,p7159,p7161,p7174,p7175);
FA fa2861(p7163,p7165,p7167,p7176,p7177);
FA fa2862(p7038,p7040,p7042,p7178,p7179);
FA fa2863(p7044,p7046,p7056,p7180,p7181);
FA fa2864(p7064,p7169,p7171,p7182,p7183);
FA fa2865(p7050,p7052,p7054,p7184,p7185);
FA fa2866(p7173,p7175,p7177,p7186,p7187);
FA fa2867(p7058,p7060,p7062,p7188,p7189);
FA fa2868(p7179,p7181,p7183,p7190,p7191);
FA fa2869(p7066,p7068,p7070,p7192,p7193);
FA fa2870(p7185,p7187,p7072,p7194,p7195);
FA fa2871(p7074,p7082,p7189,p7196,p7197);
FA fa2872(p7191,p7076,p7078,p7198,p7199);
FA fa2873(p7080,p7193,p7195,p7200,p7201);
FA fa2874(p7197,p7084,p7086,p7202,p7203);
FA fa2875(p7088,p7199,p7201,p7204,p7205);
HA ha727(p7090,p7094,p7206,p7207);
FA fa2876(p7096,p7092,p7203,p7208,p7209);
FA fa2877(p7205,p7207,p7098,p7210,p7211);
FA fa2878(p7209,p7100,p7211,p7212,p7213);
FA fa2879(p7102,p7213,p7104,p7214,p7215);
HA ha728(ip_19_63,ip_20_62,p7216,p7217);
FA fa2880(ip_21_61,ip_22_60,ip_23_59,p7218,p7219);
FA fa2881(ip_24_58,ip_25_57,ip_26_56,p7220,p7221);
FA fa2882(ip_27_55,ip_28_54,ip_29_53,p7222,p7223);
FA fa2883(ip_30_52,ip_31_51,ip_32_50,p7224,p7225);
FA fa2884(ip_33_49,ip_34_48,ip_35_47,p7226,p7227);
HA ha729(ip_36_46,ip_37_45,p7228,p7229);
FA fa2885(ip_38_44,ip_39_43,ip_40_42,p7230,p7231);
FA fa2886(ip_41_41,ip_42_40,ip_43_39,p7232,p7233);
HA ha730(ip_44_38,ip_45_37,p7234,p7235);
FA fa2887(ip_46_36,ip_47_35,ip_48_34,p7236,p7237);
FA fa2888(ip_49_33,ip_50_32,ip_51_31,p7238,p7239);
FA fa2889(ip_52_30,ip_53_29,ip_54_28,p7240,p7241);
FA fa2890(ip_55_27,ip_56_26,ip_57_25,p7242,p7243);
FA fa2891(ip_58_24,ip_59_23,ip_60_22,p7244,p7245);
HA ha731(ip_61_21,ip_62_20,p7246,p7247);
FA fa2892(ip_63_19,p7118,p7124,p7248,p7249);
FA fa2893(p7217,p7229,p7235,p7250,p7251);
FA fa2894(p7247,p7142,p7219,p7252,p7253);
FA fa2895(p7221,p7223,p7225,p7254,p7255);
FA fa2896(p7227,p7231,p7233,p7256,p7257);
FA fa2897(p7237,p7239,p7241,p7258,p7259);
FA fa2898(p7243,p7245,p7108,p7260,p7261);
FA fa2899(p7110,p7112,p7114,p7262,p7263);
FA fa2900(p7116,p7120,p7122,p7264,p7265);
FA fa2901(p7126,p7128,p7130,p7266,p7267);
FA fa2902(p7132,p7134,p7136,p7268,p7269);
FA fa2903(p7138,p7249,p7251,p7270,p7271);
FA fa2904(p7140,p7253,p7255,p7272,p7273);
FA fa2905(p7257,p7259,p7261,p7274,p7275);
FA fa2906(p7144,p7146,p7148,p7276,p7277);
FA fa2907(p7150,p7152,p7154,p7278,p7279);
FA fa2908(p7166,p7263,p7265,p7280,p7281);
FA fa2909(p7267,p7269,p7271,p7282,p7283);
HA ha732(p7156,p7158,p7284,p7285);
FA fa2910(p7160,p7162,p7164,p7286,p7287);
FA fa2911(p7273,p7275,p7168,p7288,p7289);
FA fa2912(p7170,p7277,p7279,p7290,p7291);
FA fa2913(p7281,p7283,p7285,p7292,p7293);
HA ha733(p7172,p7174,p7294,p7295);
HA ha734(p7176,p7287,p7296,p7297);
FA fa2914(p7289,p7178,p7180,p7298,p7299);
FA fa2915(p7182,p7291,p7293,p7300,p7301);
HA ha735(p7295,p7297,p7302,p7303);
FA fa2916(p7184,p7186,p7303,p7304,p7305);
FA fa2917(p7188,p7190,p7299,p7306,p7307);
FA fa2918(p7301,p7192,p7194,p7308,p7309);
FA fa2919(p7305,p7196,p7307,p7310,p7311);
FA fa2920(p7198,p7200,p7309,p7312,p7313);
HA ha736(p7206,p7311,p7314,p7315);
FA fa2921(p7202,p7204,p7313,p7316,p7317);
FA fa2922(p7315,p7208,p7317,p7318,p7319);
FA fa2923(p7210,p7319,p7212,p7320,p7321);
FA fa2924(ip_20_63,ip_21_62,ip_22_61,p7322,p7323);
FA fa2925(ip_23_60,ip_24_59,ip_25_58,p7324,p7325);
FA fa2926(ip_26_57,ip_27_56,ip_28_55,p7326,p7327);
HA ha737(ip_29_54,ip_30_53,p7328,p7329);
FA fa2927(ip_31_52,ip_32_51,ip_33_50,p7330,p7331);
FA fa2928(ip_34_49,ip_35_48,ip_36_47,p7332,p7333);
HA ha738(ip_37_46,ip_38_45,p7334,p7335);
FA fa2929(ip_39_44,ip_40_43,ip_41_42,p7336,p7337);
HA ha739(ip_42_41,ip_43_40,p7338,p7339);
FA fa2930(ip_44_39,ip_45_38,ip_46_37,p7340,p7341);
FA fa2931(ip_47_36,ip_48_35,ip_49_34,p7342,p7343);
FA fa2932(ip_50_33,ip_51_32,ip_52_31,p7344,p7345);
FA fa2933(ip_53_30,ip_54_29,ip_55_28,p7346,p7347);
FA fa2934(ip_56_27,ip_57_26,ip_58_25,p7348,p7349);
FA fa2935(ip_59_24,ip_60_23,ip_61_22,p7350,p7351);
FA fa2936(ip_62_21,ip_63_20,p7216,p7352,p7353);
HA ha740(p7228,p7234,p7354,p7355);
FA fa2937(p7246,p7329,p7335,p7356,p7357);
FA fa2938(p7339,p7323,p7325,p7358,p7359);
HA ha741(p7327,p7331,p7360,p7361);
FA fa2939(p7333,p7337,p7341,p7362,p7363);
FA fa2940(p7343,p7345,p7347,p7364,p7365);
FA fa2941(p7349,p7351,p7353,p7366,p7367);
FA fa2942(p7355,p7218,p7220,p7368,p7369);
FA fa2943(p7222,p7224,p7226,p7370,p7371);
FA fa2944(p7230,p7232,p7236,p7372,p7373);
FA fa2945(p7238,p7240,p7242,p7374,p7375);
FA fa2946(p7244,p7357,p7361,p7376,p7377);
FA fa2947(p7248,p7250,p7359,p7378,p7379);
FA fa2948(p7363,p7365,p7367,p7380,p7381);
FA fa2949(p7252,p7254,p7256,p7382,p7383);
FA fa2950(p7258,p7260,p7369,p7384,p7385);
FA fa2951(p7371,p7373,p7375,p7386,p7387);
FA fa2952(p7377,p7262,p7264,p7388,p7389);
FA fa2953(p7266,p7268,p7270,p7390,p7391);
FA fa2954(p7379,p7381,p7272,p7392,p7393);
FA fa2955(p7274,p7284,p7383,p7394,p7395);
FA fa2956(p7385,p7387,p7276,p7396,p7397);
HA ha742(p7278,p7280,p7398,p7399);
FA fa2957(p7282,p7389,p7391,p7400,p7401);
FA fa2958(p7393,p7286,p7288,p7402,p7403);
FA fa2959(p7294,p7296,p7395,p7404,p7405);
FA fa2960(p7397,p7399,p7290,p7406,p7407);
HA ha743(p7292,p7302,p7408,p7409);
HA ha744(p7401,p7403,p7410,p7411);
FA fa2961(p7405,p7407,p7409,p7412,p7413);
FA fa2962(p7298,p7300,p7411,p7414,p7415);
FA fa2963(p7304,p7413,p7306,p7416,p7417);
HA ha745(p7415,p7308,p7418,p7419);
FA fa2964(p7417,p7310,p7314,p7420,p7421);
FA fa2965(p7419,p7312,p7421,p7422,p7423);
FA fa2966(p7316,p7423,p7318,p7424,p7425);
FA fa2967(ip_21_63,ip_22_62,ip_23_61,p7426,p7427);
FA fa2968(ip_24_60,ip_25_59,ip_26_58,p7428,p7429);
FA fa2969(ip_27_57,ip_28_56,ip_29_55,p7430,p7431);
FA fa2970(ip_30_54,ip_31_53,ip_32_52,p7432,p7433);
FA fa2971(ip_33_51,ip_34_50,ip_35_49,p7434,p7435);
FA fa2972(ip_36_48,ip_37_47,ip_38_46,p7436,p7437);
FA fa2973(ip_39_45,ip_40_44,ip_41_43,p7438,p7439);
FA fa2974(ip_42_42,ip_43_41,ip_44_40,p7440,p7441);
FA fa2975(ip_45_39,ip_46_38,ip_47_37,p7442,p7443);
FA fa2976(ip_48_36,ip_49_35,ip_50_34,p7444,p7445);
FA fa2977(ip_51_33,ip_52_32,ip_53_31,p7446,p7447);
HA ha746(ip_54_30,ip_55_29,p7448,p7449);
FA fa2978(ip_56_28,ip_57_27,ip_58_26,p7450,p7451);
FA fa2979(ip_59_25,ip_60_24,ip_61_23,p7452,p7453);
FA fa2980(ip_62_22,ip_63_21,p7328,p7454,p7455);
FA fa2981(p7334,p7338,p7449,p7456,p7457);
FA fa2982(p7354,p7427,p7429,p7458,p7459);
HA ha747(p7431,p7433,p7460,p7461);
FA fa2983(p7435,p7437,p7439,p7462,p7463);
FA fa2984(p7441,p7443,p7445,p7464,p7465);
FA fa2985(p7447,p7451,p7453,p7466,p7467);
FA fa2986(p7455,p7322,p7324,p7468,p7469);
FA fa2987(p7326,p7330,p7332,p7470,p7471);
FA fa2988(p7336,p7340,p7342,p7472,p7473);
FA fa2989(p7344,p7346,p7348,p7474,p7475);
FA fa2990(p7350,p7352,p7360,p7476,p7477);
FA fa2991(p7457,p7461,p7356,p7478,p7479);
FA fa2992(p7459,p7463,p7465,p7480,p7481);
HA ha748(p7467,p7358,p7482,p7483);
FA fa2993(p7362,p7364,p7366,p7484,p7485);
FA fa2994(p7469,p7471,p7473,p7486,p7487);
FA fa2995(p7475,p7477,p7479,p7488,p7489);
FA fa2996(p7368,p7370,p7372,p7490,p7491);
FA fa2997(p7374,p7376,p7481,p7492,p7493);
FA fa2998(p7483,p7378,p7380,p7494,p7495);
FA fa2999(p7485,p7487,p7489,p7496,p7497);
FA fa3000(p7382,p7384,p7386,p7498,p7499);
FA fa3001(p7491,p7493,p7388,p7500,p7501);
HA ha749(p7390,p7392,p7502,p7503);
FA fa3002(p7398,p7495,p7497,p7504,p7505);
FA fa3003(p7394,p7396,p7499,p7506,p7507);
FA fa3004(p7501,p7503,p7400,p7508,p7509);
HA ha750(p7408,p7505,p7510,p7511);
FA fa3005(p7402,p7404,p7406,p7512,p7513);
FA fa3006(p7410,p7507,p7509,p7514,p7515);
FA fa3007(p7511,p7412,p7513,p7516,p7517);
FA fa3008(p7515,p7414,p7416,p7518,p7519);
FA fa3009(p7418,p7517,p7519,p7520,p7521);
FA fa3010(p7521,p7420,p7422,p7522,p7523);
FA fa3011(ip_22_63,ip_23_62,ip_24_61,p7524,p7525);
FA fa3012(ip_25_60,ip_26_59,ip_27_58,p7526,p7527);
FA fa3013(ip_28_57,ip_29_56,ip_30_55,p7528,p7529);
FA fa3014(ip_31_54,ip_32_53,ip_33_52,p7530,p7531);
FA fa3015(ip_34_51,ip_35_50,ip_36_49,p7532,p7533);
FA fa3016(ip_37_48,ip_38_47,ip_39_46,p7534,p7535);
FA fa3017(ip_40_45,ip_41_44,ip_42_43,p7536,p7537);
FA fa3018(ip_43_42,ip_44_41,ip_45_40,p7538,p7539);
FA fa3019(ip_46_39,ip_47_38,ip_48_37,p7540,p7541);
FA fa3020(ip_49_36,ip_50_35,ip_51_34,p7542,p7543);
HA ha751(ip_52_33,ip_53_32,p7544,p7545);
HA ha752(ip_54_31,ip_55_30,p7546,p7547);
FA fa3021(ip_56_29,ip_57_28,ip_58_27,p7548,p7549);
FA fa3022(ip_59_26,ip_60_25,ip_61_24,p7550,p7551);
HA ha753(ip_62_23,ip_63_22,p7552,p7553);
FA fa3023(p7448,p7545,p7547,p7554,p7555);
FA fa3024(p7553,p7525,p7527,p7556,p7557);
HA ha754(p7529,p7531,p7558,p7559);
HA ha755(p7533,p7535,p7560,p7561);
HA ha756(p7537,p7539,p7562,p7563);
FA fa3025(p7541,p7543,p7549,p7564,p7565);
FA fa3026(p7551,p7426,p7428,p7566,p7567);
FA fa3027(p7430,p7432,p7434,p7568,p7569);
FA fa3028(p7436,p7438,p7440,p7570,p7571);
FA fa3029(p7442,p7444,p7446,p7572,p7573);
HA ha757(p7450,p7452,p7574,p7575);
HA ha758(p7454,p7460,p7576,p7577);
FA fa3030(p7555,p7559,p7561,p7578,p7579);
FA fa3031(p7563,p7456,p7557,p7580,p7581);
HA ha759(p7565,p7575,p7582,p7583);
FA fa3032(p7577,p7458,p7462,p7584,p7585);
FA fa3033(p7464,p7466,p7567,p7586,p7587);
HA ha760(p7569,p7571,p7588,p7589);
FA fa3034(p7573,p7579,p7583,p7590,p7591);
FA fa3035(p7468,p7470,p7472,p7592,p7593);
FA fa3036(p7474,p7476,p7478,p7594,p7595);
FA fa3037(p7482,p7581,p7589,p7596,p7597);
FA fa3038(p7480,p7585,p7587,p7598,p7599);
FA fa3039(p7591,p7484,p7486,p7600,p7601);
FA fa3040(p7488,p7593,p7595,p7602,p7603);
FA fa3041(p7597,p7490,p7492,p7604,p7605);
FA fa3042(p7599,p7494,p7496,p7606,p7607);
FA fa3043(p7502,p7601,p7603,p7608,p7609);
FA fa3044(p7498,p7500,p7605,p7610,p7611);
FA fa3045(p7504,p7510,p7607,p7612,p7613);
FA fa3046(p7609,p7506,p7508,p7614,p7615);
FA fa3047(p7611,p7613,p7512,p7616,p7617);
FA fa3048(p7514,p7615,p7617,p7618,p7619);
FA fa3049(p7516,p7619,p7518,p7620,p7621);
HA ha761(p7520,p7621,p7622,p7623);
FA fa3050(ip_23_63,ip_24_62,ip_25_61,p7624,p7625);
HA ha762(ip_26_60,ip_27_59,p7626,p7627);
FA fa3051(ip_28_58,ip_29_57,ip_30_56,p7628,p7629);
FA fa3052(ip_31_55,ip_32_54,ip_33_53,p7630,p7631);
HA ha763(ip_34_52,ip_35_51,p7632,p7633);
FA fa3053(ip_36_50,ip_37_49,ip_38_48,p7634,p7635);
FA fa3054(ip_39_47,ip_40_46,ip_41_45,p7636,p7637);
FA fa3055(ip_42_44,ip_43_43,ip_44_42,p7638,p7639);
FA fa3056(ip_45_41,ip_46_40,ip_47_39,p7640,p7641);
FA fa3057(ip_48_38,ip_49_37,ip_50_36,p7642,p7643);
FA fa3058(ip_51_35,ip_52_34,ip_53_33,p7644,p7645);
FA fa3059(ip_54_32,ip_55_31,ip_56_30,p7646,p7647);
FA fa3060(ip_57_29,ip_58_28,ip_59_27,p7648,p7649);
HA ha764(ip_60_26,ip_61_25,p7650,p7651);
FA fa3061(ip_62_24,ip_63_23,p7544,p7652,p7653);
FA fa3062(p7546,p7552,p7627,p7654,p7655);
FA fa3063(p7633,p7651,p7625,p7656,p7657);
FA fa3064(p7629,p7631,p7635,p7658,p7659);
FA fa3065(p7637,p7639,p7641,p7660,p7661);
FA fa3066(p7643,p7645,p7647,p7662,p7663);
FA fa3067(p7649,p7653,p7524,p7664,p7665);
FA fa3068(p7526,p7528,p7530,p7666,p7667);
HA ha765(p7532,p7534,p7668,p7669);
FA fa3069(p7536,p7538,p7540,p7670,p7671);
HA ha766(p7542,p7548,p7672,p7673);
FA fa3070(p7550,p7558,p7560,p7674,p7675);
FA fa3071(p7562,p7655,p7657,p7676,p7677);
FA fa3072(p7554,p7574,p7576,p7678,p7679);
FA fa3073(p7659,p7661,p7663,p7680,p7681);
HA ha767(p7665,p7669,p7682,p7683);
FA fa3074(p7673,p7556,p7564,p7684,p7685);
FA fa3075(p7582,p7667,p7671,p7686,p7687);
FA fa3076(p7675,p7677,p7683,p7688,p7689);
HA ha768(p7566,p7568,p7690,p7691);
FA fa3077(p7570,p7572,p7578,p7692,p7693);
FA fa3078(p7588,p7679,p7681,p7694,p7695);
FA fa3079(p7580,p7685,p7687,p7696,p7697);
FA fa3080(p7689,p7691,p7584,p7698,p7699);
FA fa3081(p7586,p7590,p7693,p7700,p7701);
FA fa3082(p7695,p7592,p7594,p7702,p7703);
FA fa3083(p7596,p7697,p7699,p7704,p7705);
FA fa3084(p7598,p7701,p7600,p7706,p7707);
FA fa3085(p7602,p7703,p7705,p7708,p7709);
FA fa3086(p7604,p7707,p7606,p7710,p7711);
FA fa3087(p7608,p7709,p7610,p7712,p7713);
FA fa3088(p7711,p7612,p7713,p7714,p7715);
FA fa3089(p7614,p7616,p7715,p7716,p7717);
FA fa3090(p7618,p7717,p7620,p7718,p7719);
FA fa3091(ip_24_63,ip_25_62,ip_26_61,p7720,p7721);
FA fa3092(ip_27_60,ip_28_59,ip_29_58,p7722,p7723);
FA fa3093(ip_30_57,ip_31_56,ip_32_55,p7724,p7725);
FA fa3094(ip_33_54,ip_34_53,ip_35_52,p7726,p7727);
FA fa3095(ip_36_51,ip_37_50,ip_38_49,p7728,p7729);
HA ha769(ip_39_48,ip_40_47,p7730,p7731);
FA fa3096(ip_41_46,ip_42_45,ip_43_44,p7732,p7733);
FA fa3097(ip_44_43,ip_45_42,ip_46_41,p7734,p7735);
HA ha770(ip_47_40,ip_48_39,p7736,p7737);
FA fa3098(ip_49_38,ip_50_37,ip_51_36,p7738,p7739);
FA fa3099(ip_52_35,ip_53_34,ip_54_33,p7740,p7741);
FA fa3100(ip_55_32,ip_56_31,ip_57_30,p7742,p7743);
FA fa3101(ip_58_29,ip_59_28,ip_60_27,p7744,p7745);
FA fa3102(ip_61_26,ip_62_25,ip_63_24,p7746,p7747);
FA fa3103(p7626,p7632,p7650,p7748,p7749);
FA fa3104(p7731,p7737,p7721,p7750,p7751);
FA fa3105(p7723,p7725,p7727,p7752,p7753);
FA fa3106(p7729,p7733,p7735,p7754,p7755);
FA fa3107(p7739,p7741,p7743,p7756,p7757);
FA fa3108(p7745,p7747,p7624,p7758,p7759);
FA fa3109(p7628,p7630,p7634,p7760,p7761);
FA fa3110(p7636,p7638,p7640,p7762,p7763);
FA fa3111(p7642,p7644,p7646,p7764,p7765);
HA ha771(p7648,p7652,p7766,p7767);
HA ha772(p7749,p7751,p7768,p7769);
FA fa3112(p7654,p7656,p7668,p7770,p7771);
FA fa3113(p7672,p7753,p7755,p7772,p7773);
FA fa3114(p7757,p7759,p7767,p7774,p7775);
FA fa3115(p7769,p7658,p7660,p7776,p7777);
FA fa3116(p7662,p7664,p7682,p7778,p7779);
FA fa3117(p7761,p7763,p7765,p7780,p7781);
FA fa3118(p7666,p7670,p7674,p7782,p7783);
FA fa3119(p7676,p7771,p7773,p7784,p7785);
FA fa3120(p7775,p7678,p7680,p7786,p7787);
FA fa3121(p7690,p7777,p7779,p7788,p7789);
FA fa3122(p7781,p7684,p7686,p7790,p7791);
FA fa3123(p7688,p7783,p7785,p7792,p7793);
FA fa3124(p7692,p7694,p7787,p7794,p7795);
FA fa3125(p7789,p7696,p7698,p7796,p7797);
FA fa3126(p7791,p7793,p7700,p7798,p7799);
FA fa3127(p7795,p7702,p7704,p7800,p7801);
FA fa3128(p7797,p7799,p7706,p7802,p7803);
FA fa3129(p7708,p7801,p7803,p7804,p7805);
FA fa3130(p7710,p7712,p7805,p7806,p7807);
FA fa3131(p7714,p7807,p7716,p7808,p7809);
HA ha773(ip_25_63,ip_26_62,p7810,p7811);
FA fa3132(ip_27_61,ip_28_60,ip_29_59,p7812,p7813);
FA fa3133(ip_30_58,ip_31_57,ip_32_56,p7814,p7815);
FA fa3134(ip_33_55,ip_34_54,ip_35_53,p7816,p7817);
HA ha774(ip_36_52,ip_37_51,p7818,p7819);
HA ha775(ip_38_50,ip_39_49,p7820,p7821);
FA fa3135(ip_40_48,ip_41_47,ip_42_46,p7822,p7823);
FA fa3136(ip_43_45,ip_44_44,ip_45_43,p7824,p7825);
HA ha776(ip_46_42,ip_47_41,p7826,p7827);
FA fa3137(ip_48_40,ip_49_39,ip_50_38,p7828,p7829);
FA fa3138(ip_51_37,ip_52_36,ip_53_35,p7830,p7831);
FA fa3139(ip_54_34,ip_55_33,ip_56_32,p7832,p7833);
FA fa3140(ip_57_31,ip_58_30,ip_59_29,p7834,p7835);
FA fa3141(ip_60_28,ip_61_27,ip_62_26,p7836,p7837);
FA fa3142(ip_63_25,p7730,p7736,p7838,p7839);
HA ha777(p7811,p7819,p7840,p7841);
FA fa3143(p7821,p7827,p7813,p7842,p7843);
FA fa3144(p7815,p7817,p7823,p7844,p7845);
FA fa3145(p7825,p7829,p7831,p7846,p7847);
FA fa3146(p7833,p7835,p7837,p7848,p7849);
FA fa3147(p7841,p7720,p7722,p7850,p7851);
HA ha778(p7724,p7726,p7852,p7853);
HA ha779(p7728,p7732,p7854,p7855);
FA fa3148(p7734,p7738,p7740,p7856,p7857);
FA fa3149(p7742,p7744,p7746,p7858,p7859);
HA ha780(p7839,p7843,p7860,p7861);
FA fa3150(p7748,p7750,p7766,p7862,p7863);
FA fa3151(p7768,p7845,p7847,p7864,p7865);
FA fa3152(p7849,p7853,p7855,p7866,p7867);
FA fa3153(p7861,p7752,p7754,p7868,p7869);
FA fa3154(p7756,p7758,p7851,p7870,p7871);
FA fa3155(p7857,p7859,p7760,p7872,p7873);
HA ha781(p7762,p7764,p7874,p7875);
FA fa3156(p7863,p7865,p7867,p7876,p7877);
FA fa3157(p7770,p7772,p7774,p7878,p7879);
FA fa3158(p7869,p7871,p7873,p7880,p7881);
FA fa3159(p7875,p7776,p7778,p7882,p7883);
FA fa3160(p7780,p7877,p7782,p7884,p7885);
FA fa3161(p7784,p7879,p7881,p7886,p7887);
FA fa3162(p7786,p7788,p7883,p7888,p7889);
FA fa3163(p7885,p7790,p7792,p7890,p7891);
FA fa3164(p7887,p7794,p7889,p7892,p7893);
FA fa3165(p7796,p7798,p7891,p7894,p7895);
FA fa3166(p7893,p7800,p7802,p7896,p7897);
FA fa3167(p7895,p7804,p7897,p7898,p7899);
FA fa3168(p7806,p7899,p7808,p7900,p7901);
FA fa3169(ip_26_63,ip_27_62,ip_28_61,p7902,p7903);
FA fa3170(ip_29_60,ip_30_59,ip_31_58,p7904,p7905);
HA ha782(ip_32_57,ip_33_56,p7906,p7907);
FA fa3171(ip_34_55,ip_35_54,ip_36_53,p7908,p7909);
FA fa3172(ip_37_52,ip_38_51,ip_39_50,p7910,p7911);
FA fa3173(ip_40_49,ip_41_48,ip_42_47,p7912,p7913);
HA ha783(ip_43_46,ip_44_45,p7914,p7915);
FA fa3174(ip_45_44,ip_46_43,ip_47_42,p7916,p7917);
FA fa3175(ip_48_41,ip_49_40,ip_50_39,p7918,p7919);
FA fa3176(ip_51_38,ip_52_37,ip_53_36,p7920,p7921);
FA fa3177(ip_54_35,ip_55_34,ip_56_33,p7922,p7923);
FA fa3178(ip_57_32,ip_58_31,ip_59_30,p7924,p7925);
HA ha784(ip_60_29,ip_61_28,p7926,p7927);
FA fa3179(ip_62_27,ip_63_26,p7810,p7928,p7929);
FA fa3180(p7818,p7820,p7826,p7930,p7931);
HA ha785(p7907,p7915,p7932,p7933);
FA fa3181(p7927,p7840,p7903,p7934,p7935);
FA fa3182(p7905,p7909,p7911,p7936,p7937);
FA fa3183(p7913,p7917,p7919,p7938,p7939);
HA ha786(p7921,p7923,p7940,p7941);
FA fa3184(p7925,p7929,p7933,p7942,p7943);
FA fa3185(p7812,p7814,p7816,p7944,p7945);
FA fa3186(p7822,p7824,p7828,p7946,p7947);
FA fa3187(p7830,p7832,p7834,p7948,p7949);
FA fa3188(p7836,p7931,p7941,p7950,p7951);
FA fa3189(p7838,p7842,p7852,p7952,p7953);
FA fa3190(p7854,p7860,p7935,p7954,p7955);
FA fa3191(p7937,p7939,p7943,p7956,p7957);
FA fa3192(p7844,p7846,p7848,p7958,p7959);
HA ha787(p7945,p7947,p7960,p7961);
FA fa3193(p7949,p7951,p7850,p7962,p7963);
FA fa3194(p7856,p7858,p7953,p7964,p7965);
FA fa3195(p7955,p7957,p7961,p7966,p7967);
HA ha788(p7862,p7864,p7968,p7969);
FA fa3196(p7866,p7874,p7959,p7970,p7971);
FA fa3197(p7963,p7868,p7870,p7972,p7973);
FA fa3198(p7872,p7965,p7967,p7974,p7975);
FA fa3199(p7969,p7876,p7971,p7976,p7977);
FA fa3200(p7878,p7880,p7973,p7978,p7979);
FA fa3201(p7975,p7882,p7884,p7980,p7981);
FA fa3202(p7977,p7886,p7979,p7982,p7983);
FA fa3203(p7888,p7981,p7890,p7984,p7985);
FA fa3204(p7983,p7892,p7985,p7986,p7987);
FA fa3205(p7894,p7987,p7896,p7988,p7989);
FA fa3206(p7989,p7898,p7900,p7990,p7991);
FA fa3207(ip_27_63,ip_28_62,ip_29_61,p7992,p7993);
FA fa3208(ip_30_60,ip_31_59,ip_32_58,p7994,p7995);
FA fa3209(ip_33_57,ip_34_56,ip_35_55,p7996,p7997);
FA fa3210(ip_36_54,ip_37_53,ip_38_52,p7998,p7999);
FA fa3211(ip_39_51,ip_40_50,ip_41_49,p8000,p8001);
FA fa3212(ip_42_48,ip_43_47,ip_44_46,p8002,p8003);
FA fa3213(ip_45_45,ip_46_44,ip_47_43,p8004,p8005);
FA fa3214(ip_48_42,ip_49_41,ip_50_40,p8006,p8007);
FA fa3215(ip_51_39,ip_52_38,ip_53_37,p8008,p8009);
HA ha789(ip_54_36,ip_55_35,p8010,p8011);
FA fa3216(ip_56_34,ip_57_33,ip_58_32,p8012,p8013);
FA fa3217(ip_59_31,ip_60_30,ip_61_29,p8014,p8015);
FA fa3218(ip_62_28,ip_63_27,p7906,p8016,p8017);
FA fa3219(p7914,p7926,p8011,p8018,p8019);
HA ha790(p7932,p7993,p8020,p8021);
FA fa3220(p7995,p7997,p7999,p8022,p8023);
FA fa3221(p8001,p8003,p8005,p8024,p8025);
FA fa3222(p8007,p8009,p8013,p8026,p8027);
FA fa3223(p8015,p8017,p7902,p8028,p8029);
FA fa3224(p7904,p7908,p7910,p8030,p8031);
FA fa3225(p7912,p7916,p7918,p8032,p8033);
FA fa3226(p7920,p7922,p7924,p8034,p8035);
FA fa3227(p7928,p7940,p8019,p8036,p8037);
FA fa3228(p8021,p7930,p8023,p8038,p8039);
FA fa3229(p8025,p8027,p8029,p8040,p8041);
FA fa3230(p7934,p7936,p7938,p8042,p8043);
FA fa3231(p7942,p8031,p8033,p8044,p8045);
FA fa3232(p8035,p8037,p7944,p8046,p8047);
HA ha791(p7946,p7948,p8048,p8049);
FA fa3233(p7950,p7960,p8039,p8050,p8051);
FA fa3234(p8041,p7952,p7954,p8052,p8053);
HA ha792(p7956,p8043,p8054,p8055);
FA fa3235(p8045,p8047,p8049,p8056,p8057);
FA fa3236(p7958,p7962,p7968,p8058,p8059);
FA fa3237(p8051,p8055,p7964,p8060,p8061);
FA fa3238(p7966,p8053,p8057,p8062,p8063);
FA fa3239(p7970,p8059,p8061,p8064,p8065);
FA fa3240(p7972,p7974,p8063,p8066,p8067);
FA fa3241(p7976,p8065,p7978,p8068,p8069);
FA fa3242(p8067,p7980,p8069,p8070,p8071);
HA ha793(p7982,p7984,p8072,p8073);
HA ha794(p8071,p8073,p8074,p8075);
FA fa3243(p7986,p8075,p7988,p8076,p8077);
FA fa3244(ip_28_63,ip_29_62,ip_30_61,p8078,p8079);
FA fa3245(ip_31_60,ip_32_59,ip_33_58,p8080,p8081);
FA fa3246(ip_34_57,ip_35_56,ip_36_55,p8082,p8083);
HA ha795(ip_37_54,ip_38_53,p8084,p8085);
FA fa3247(ip_39_52,ip_40_51,ip_41_50,p8086,p8087);
FA fa3248(ip_42_49,ip_43_48,ip_44_47,p8088,p8089);
HA ha796(ip_45_46,ip_46_45,p8090,p8091);
HA ha797(ip_47_44,ip_48_43,p8092,p8093);
FA fa3249(ip_49_42,ip_50_41,ip_51_40,p8094,p8095);
HA ha798(ip_52_39,ip_53_38,p8096,p8097);
FA fa3250(ip_54_37,ip_55_36,ip_56_35,p8098,p8099);
FA fa3251(ip_57_34,ip_58_33,ip_59_32,p8100,p8101);
FA fa3252(ip_60_31,ip_61_30,ip_62_29,p8102,p8103);
FA fa3253(ip_63_28,p8010,p8085,p8104,p8105);
FA fa3254(p8091,p8093,p8097,p8106,p8107);
FA fa3255(p8079,p8081,p8083,p8108,p8109);
HA ha799(p8087,p8089,p8110,p8111);
FA fa3256(p8095,p8099,p8101,p8112,p8113);
HA ha800(p8103,p7992,p8114,p8115);
FA fa3257(p7994,p7996,p7998,p8116,p8117);
FA fa3258(p8000,p8002,p8004,p8118,p8119);
HA ha801(p8006,p8008,p8120,p8121);
FA fa3259(p8012,p8014,p8016,p8122,p8123);
HA ha802(p8020,p8105,p8124,p8125);
FA fa3260(p8107,p8111,p8018,p8126,p8127);
HA ha803(p8109,p8113,p8128,p8129);
FA fa3261(p8115,p8121,p8125,p8130,p8131);
HA ha804(p8022,p8024,p8132,p8133);
FA fa3262(p8026,p8028,p8117,p8134,p8135);
FA fa3263(p8119,p8123,p8127,p8136,p8137);
FA fa3264(p8129,p8030,p8032,p8138,p8139);
FA fa3265(p8034,p8036,p8131,p8140,p8141);
FA fa3266(p8133,p8038,p8040,p8142,p8143);
FA fa3267(p8048,p8135,p8137,p8144,p8145);
FA fa3268(p8042,p8044,p8046,p8146,p8147);
FA fa3269(p8054,p8139,p8141,p8148,p8149);
FA fa3270(p8050,p8143,p8145,p8150,p8151);
FA fa3271(p8052,p8056,p8147,p8152,p8153);
FA fa3272(p8149,p8058,p8060,p8154,p8155);
FA fa3273(p8151,p8062,p8153,p8156,p8157);
FA fa3274(p8064,p8155,p8066,p8158,p8159);
FA fa3275(p8157,p8068,p8159,p8160,p8161);
FA fa3276(p8070,p8072,p8161,p8162,p8163);
HA ha805(p8074,p8163,p8164,p8165);
FA fa3277(ip_29_63,ip_30_62,ip_31_61,p8166,p8167);
FA fa3278(ip_32_60,ip_33_59,ip_34_58,p8168,p8169);
FA fa3279(ip_35_57,ip_36_56,ip_37_55,p8170,p8171);
FA fa3280(ip_38_54,ip_39_53,ip_40_52,p8172,p8173);
FA fa3281(ip_41_51,ip_42_50,ip_43_49,p8174,p8175);
HA ha806(ip_44_48,ip_45_47,p8176,p8177);
FA fa3282(ip_46_46,ip_47_45,ip_48_44,p8178,p8179);
FA fa3283(ip_49_43,ip_50_42,ip_51_41,p8180,p8181);
HA ha807(ip_52_40,ip_53_39,p8182,p8183);
FA fa3284(ip_54_38,ip_55_37,ip_56_36,p8184,p8185);
FA fa3285(ip_57_35,ip_58_34,ip_59_33,p8186,p8187);
FA fa3286(ip_60_32,ip_61_31,ip_62_30,p8188,p8189);
FA fa3287(ip_63_29,p8084,p8090,p8190,p8191);
FA fa3288(p8092,p8096,p8177,p8192,p8193);
FA fa3289(p8183,p8167,p8169,p8194,p8195);
HA ha808(p8171,p8173,p8196,p8197);
FA fa3290(p8175,p8179,p8181,p8198,p8199);
FA fa3291(p8185,p8187,p8189,p8200,p8201);
FA fa3292(p8078,p8080,p8082,p8202,p8203);
FA fa3293(p8086,p8088,p8094,p8204,p8205);
FA fa3294(p8098,p8100,p8102,p8206,p8207);
FA fa3295(p8110,p8191,p8193,p8208,p8209);
FA fa3296(p8197,p8104,p8106,p8210,p8211);
FA fa3297(p8114,p8120,p8124,p8212,p8213);
FA fa3298(p8195,p8199,p8201,p8214,p8215);
FA fa3299(p8108,p8112,p8128,p8216,p8217);
FA fa3300(p8203,p8205,p8207,p8218,p8219);
FA fa3301(p8209,p8116,p8118,p8220,p8221);
HA ha809(p8122,p8126,p8222,p8223);
FA fa3302(p8132,p8211,p8213,p8224,p8225);
FA fa3303(p8215,p8130,p8217,p8226,p8227);
FA fa3304(p8219,p8223,p8134,p8228,p8229);
FA fa3305(p8136,p8221,p8225,p8230,p8231);
FA fa3306(p8138,p8140,p8227,p8232,p8233);
HA ha810(p8229,p8142,p8234,p8235);
FA fa3307(p8144,p8231,p8146,p8236,p8237);
FA fa3308(p8148,p8233,p8235,p8238,p8239);
HA ha811(p8150,p8237,p8240,p8241);
FA fa3309(p8152,p8239,p8241,p8242,p8243);
FA fa3310(p8154,p8156,p8243,p8244,p8245);
FA fa3311(p8158,p8245,p8160,p8246,p8247);
FA fa3312(p8247,p8162,p8164,p8248,p8249);
FA fa3313(ip_30_63,ip_31_62,ip_32_61,p8250,p8251);
FA fa3314(ip_33_60,ip_34_59,ip_35_58,p8252,p8253);
FA fa3315(ip_36_57,ip_37_56,ip_38_55,p8254,p8255);
FA fa3316(ip_39_54,ip_40_53,ip_41_52,p8256,p8257);
FA fa3317(ip_42_51,ip_43_50,ip_44_49,p8258,p8259);
FA fa3318(ip_45_48,ip_46_47,ip_47_46,p8260,p8261);
FA fa3319(ip_48_45,ip_49_44,ip_50_43,p8262,p8263);
FA fa3320(ip_51_42,ip_52_41,ip_53_40,p8264,p8265);
HA ha812(ip_54_39,ip_55_38,p8266,p8267);
FA fa3321(ip_56_37,ip_57_36,ip_58_35,p8268,p8269);
FA fa3322(ip_59_34,ip_60_33,ip_61_32,p8270,p8271);
FA fa3323(ip_62_31,ip_63_30,p8176,p8272,p8273);
FA fa3324(p8182,p8267,p8251,p8274,p8275);
FA fa3325(p8253,p8255,p8257,p8276,p8277);
FA fa3326(p8259,p8261,p8263,p8278,p8279);
FA fa3327(p8265,p8269,p8271,p8280,p8281);
FA fa3328(p8273,p8166,p8168,p8282,p8283);
FA fa3329(p8170,p8172,p8174,p8284,p8285);
FA fa3330(p8178,p8180,p8184,p8286,p8287);
FA fa3331(p8186,p8188,p8196,p8288,p8289);
FA fa3332(p8275,p8190,p8192,p8290,p8291);
FA fa3333(p8277,p8279,p8281,p8292,p8293);
HA ha813(p8194,p8198,p8294,p8295);
HA ha814(p8200,p8283,p8296,p8297);
HA ha815(p8285,p8287,p8298,p8299);
HA ha816(p8289,p8202,p8300,p8301);
FA fa3334(p8204,p8206,p8208,p8302,p8303);
HA ha817(p8291,p8293,p8304,p8305);
FA fa3335(p8295,p8297,p8299,p8306,p8307);
FA fa3336(p8210,p8212,p8214,p8308,p8309);
FA fa3337(p8222,p8301,p8305,p8310,p8311);
HA ha818(p8216,p8218,p8312,p8313);
HA ha819(p8303,p8307,p8314,p8315);
HA ha820(p8220,p8224,p8316,p8317);
FA fa3338(p8309,p8311,p8313,p8318,p8319);
FA fa3339(p8315,p8226,p8228,p8320,p8321);
HA ha821(p8317,p8230,p8322,p8323);
FA fa3340(p8234,p8319,p8232,p8324,p8325);
HA ha822(p8321,p8323,p8326,p8327);
FA fa3341(p8236,p8240,p8325,p8328,p8329);
FA fa3342(p8327,p8238,p8329,p8330,p8331);
FA fa3343(p8242,p8331,p8244,p8332,p8333);
FA fa3344(p8333,p8246,p8248,p8334,p8335);
FA fa3345(ip_31_63,ip_32_62,ip_33_61,p8336,p8337);
FA fa3346(ip_34_60,ip_35_59,ip_36_58,p8338,p8339);
FA fa3347(ip_37_57,ip_38_56,ip_39_55,p8340,p8341);
FA fa3348(ip_40_54,ip_41_53,ip_42_52,p8342,p8343);
FA fa3349(ip_43_51,ip_44_50,ip_45_49,p8344,p8345);
FA fa3350(ip_46_48,ip_47_47,ip_48_46,p8346,p8347);
FA fa3351(ip_49_45,ip_50_44,ip_51_43,p8348,p8349);
FA fa3352(ip_52_42,ip_53_41,ip_54_40,p8350,p8351);
FA fa3353(ip_55_39,ip_56_38,ip_57_37,p8352,p8353);
FA fa3354(ip_58_36,ip_59_35,ip_60_34,p8354,p8355);
HA ha823(ip_61_33,ip_62_32,p8356,p8357);
FA fa3355(ip_63_31,p8266,p8357,p8358,p8359);
FA fa3356(p8337,p8339,p8341,p8360,p8361);
FA fa3357(p8343,p8345,p8347,p8362,p8363);
FA fa3358(p8349,p8351,p8353,p8364,p8365);
FA fa3359(p8355,p8250,p8252,p8366,p8367);
FA fa3360(p8254,p8256,p8258,p8368,p8369);
FA fa3361(p8260,p8262,p8264,p8370,p8371);
FA fa3362(p8268,p8270,p8272,p8372,p8373);
FA fa3363(p8359,p8274,p8361,p8374,p8375);
FA fa3364(p8363,p8365,p8276,p8376,p8377);
FA fa3365(p8278,p8280,p8367,p8378,p8379);
FA fa3366(p8369,p8371,p8373,p8380,p8381);
FA fa3367(p8282,p8284,p8286,p8382,p8383);
FA fa3368(p8288,p8294,p8296,p8384,p8385);
FA fa3369(p8298,p8375,p8377,p8386,p8387);
HA ha824(p8290,p8292,p8388,p8389);
FA fa3370(p8300,p8304,p8379,p8390,p8391);
HA ha825(p8381,p8383,p8392,p8393);
FA fa3371(p8385,p8387,p8389,p8394,p8395);
FA fa3372(p8302,p8306,p8312,p8396,p8397);
FA fa3373(p8314,p8391,p8393,p8398,p8399);
FA fa3374(p8308,p8310,p8316,p8400,p8401);
FA fa3375(p8395,p8397,p8399,p8402,p8403);
FA fa3376(p8318,p8322,p8401,p8404,p8405);
FA fa3377(p8320,p8326,p8403,p8406,p8407);
HA ha826(p8324,p8405,p8408,p8409);
FA fa3378(p8407,p8409,p8328,p8410,p8411);
FA fa3379(p8330,p8411,p8332,p8412,p8413);
FA fa3380(ip_32_63,ip_33_62,ip_34_61,p8414,p8415);
FA fa3381(ip_35_60,ip_36_59,ip_37_58,p8416,p8417);
FA fa3382(ip_38_57,ip_39_56,ip_40_55,p8418,p8419);
FA fa3383(ip_41_54,ip_42_53,ip_43_52,p8420,p8421);
FA fa3384(ip_44_51,ip_45_50,ip_46_49,p8422,p8423);
FA fa3385(ip_47_48,ip_48_47,ip_49_46,p8424,p8425);
FA fa3386(ip_50_45,ip_51_44,ip_52_43,p8426,p8427);
FA fa3387(ip_53_42,ip_54_41,ip_55_40,p8428,p8429);
FA fa3388(ip_56_39,ip_57_38,ip_58_37,p8430,p8431);
FA fa3389(ip_59_36,ip_60_35,ip_61_34,p8432,p8433);
FA fa3390(ip_62_33,ip_63_32,p8356,p8434,p8435);
FA fa3391(p8415,p8417,p8419,p8436,p8437);
FA fa3392(p8421,p8423,p8425,p8438,p8439);
HA ha827(p8427,p8429,p8440,p8441);
FA fa3393(p8431,p8433,p8435,p8442,p8443);
FA fa3394(p8336,p8338,p8340,p8444,p8445);
FA fa3395(p8342,p8344,p8346,p8446,p8447);
FA fa3396(p8348,p8350,p8352,p8448,p8449);
FA fa3397(p8354,p8441,p8358,p8450,p8451);
FA fa3398(p8437,p8439,p8443,p8452,p8453);
FA fa3399(p8360,p8362,p8364,p8454,p8455);
HA ha828(p8445,p8447,p8456,p8457);
HA ha829(p8449,p8451,p8458,p8459);
FA fa3400(p8366,p8368,p8370,p8460,p8461);
FA fa3401(p8372,p8453,p8457,p8462,p8463);
FA fa3402(p8459,p8374,p8376,p8464,p8465);
HA ha830(p8455,p8378,p8466,p8467);
FA fa3403(p8380,p8388,p8461,p8468,p8469);
FA fa3404(p8463,p8382,p8384,p8470,p8471);
FA fa3405(p8386,p8392,p8465,p8472,p8473);
HA ha831(p8467,p8390,p8474,p8475);
HA ha832(p8469,p8394,p8476,p8477);
FA fa3406(p8471,p8473,p8475,p8478,p8479);
HA ha833(p8396,p8398,p8480,p8481);
HA ha834(p8477,p8400,p8482,p8483);
FA fa3407(p8479,p8481,p8402,p8484,p8485);
FA fa3408(p8483,p8404,p8408,p8486,p8487);
FA fa3409(p8485,p8406,p8487,p8488,p8489);
FA fa3410(p8410,p8489,p8412,p8490,p8491);
FA fa3411(ip_33_63,ip_34_62,ip_35_61,p8492,p8493);
FA fa3412(ip_36_60,ip_37_59,ip_38_58,p8494,p8495);
HA ha835(ip_39_57,ip_40_56,p8496,p8497);
FA fa3413(ip_41_55,ip_42_54,ip_43_53,p8498,p8499);
FA fa3414(ip_44_52,ip_45_51,ip_46_50,p8500,p8501);
FA fa3415(ip_47_49,ip_48_48,ip_49_47,p8502,p8503);
FA fa3416(ip_50_46,ip_51_45,ip_52_44,p8504,p8505);
HA ha836(ip_53_43,ip_54_42,p8506,p8507);
FA fa3417(ip_55_41,ip_56_40,ip_57_39,p8508,p8509);
FA fa3418(ip_58_38,ip_59_37,ip_60_36,p8510,p8511);
FA fa3419(ip_61_35,ip_62_34,ip_63_33,p8512,p8513);
HA ha837(p8497,p8507,p8514,p8515);
FA fa3420(p8493,p8495,p8499,p8516,p8517);
FA fa3421(p8501,p8503,p8505,p8518,p8519);
FA fa3422(p8509,p8511,p8513,p8520,p8521);
FA fa3423(p8515,p8414,p8416,p8522,p8523);
FA fa3424(p8418,p8420,p8422,p8524,p8525);
FA fa3425(p8424,p8426,p8428,p8526,p8527);
FA fa3426(p8430,p8432,p8434,p8528,p8529);
FA fa3427(p8440,p8517,p8519,p8530,p8531);
FA fa3428(p8521,p8436,p8438,p8532,p8533);
FA fa3429(p8442,p8523,p8525,p8534,p8535);
FA fa3430(p8527,p8529,p8444,p8536,p8537);
FA fa3431(p8446,p8448,p8450,p8538,p8539);
FA fa3432(p8456,p8458,p8531,p8540,p8541);
FA fa3433(p8452,p8533,p8535,p8542,p8543);
FA fa3434(p8537,p8454,p8539,p8544,p8545);
FA fa3435(p8541,p8460,p8462,p8546,p8547);
FA fa3436(p8466,p8543,p8464,p8548,p8549);
FA fa3437(p8545,p8468,p8474,p8550,p8551);
FA fa3438(p8547,p8549,p8470,p8552,p8553);
FA fa3439(p8472,p8476,p8480,p8554,p8555);
FA fa3440(p8551,p8553,p8478,p8556,p8557);
FA fa3441(p8482,p8555,p8557,p8558,p8559);
HA ha838(p8484,p8559,p8560,p8561);
FA fa3442(p8561,p8486,p8488,p8562,p8563);
HA ha839(ip_34_63,ip_35_62,p8564,p8565);
FA fa3443(ip_36_61,ip_37_60,ip_38_59,p8566,p8567);
FA fa3444(ip_39_58,ip_40_57,ip_41_56,p8568,p8569);
FA fa3445(ip_42_55,ip_43_54,ip_44_53,p8570,p8571);
FA fa3446(ip_45_52,ip_46_51,ip_47_50,p8572,p8573);
HA ha840(ip_48_49,ip_49_48,p8574,p8575);
HA ha841(ip_50_47,ip_51_46,p8576,p8577);
FA fa3447(ip_52_45,ip_53_44,ip_54_43,p8578,p8579);
FA fa3448(ip_55_42,ip_56_41,ip_57_40,p8580,p8581);
FA fa3449(ip_58_39,ip_59_38,ip_60_37,p8582,p8583);
FA fa3450(ip_61_36,ip_62_35,ip_63_34,p8584,p8585);
FA fa3451(p8496,p8506,p8565,p8586,p8587);
FA fa3452(p8575,p8577,p8514,p8588,p8589);
FA fa3453(p8567,p8569,p8571,p8590,p8591);
FA fa3454(p8573,p8579,p8581,p8592,p8593);
FA fa3455(p8583,p8585,p8492,p8594,p8595);
HA ha842(p8494,p8498,p8596,p8597);
FA fa3456(p8500,p8502,p8504,p8598,p8599);
FA fa3457(p8508,p8510,p8512,p8600,p8601);
FA fa3458(p8587,p8589,p8591,p8602,p8603);
HA ha843(p8593,p8595,p8604,p8605);
FA fa3459(p8597,p8516,p8518,p8606,p8607);
FA fa3460(p8520,p8599,p8601,p8608,p8609);
FA fa3461(p8603,p8605,p8522,p8610,p8611);
FA fa3462(p8524,p8526,p8528,p8612,p8613);
FA fa3463(p8530,p8607,p8609,p8614,p8615);
HA ha844(p8611,p8532,p8616,p8617);
FA fa3464(p8534,p8536,p8613,p8618,p8619);
FA fa3465(p8538,p8540,p8615,p8620,p8621);
FA fa3466(p8617,p8542,p8619,p8622,p8623);
HA ha845(p8544,p8621,p8624,p8625);
HA ha846(p8546,p8548,p8626,p8627);
HA ha847(p8623,p8625,p8628,p8629);
HA ha848(p8627,p8629,p8630,p8631);
HA ha849(p8550,p8552,p8632,p8633);
HA ha850(p8631,p8554,p8634,p8635);
HA ha851(p8633,p8556,p8636,p8637);
FA fa3467(p8635,p8558,p8560,p8638,p8639);
FA fa3468(p8637,p8639,p8562,p8640,p8641);
FA fa3469(ip_35_63,ip_36_62,ip_37_61,p8642,p8643);
HA ha852(ip_38_60,ip_39_59,p8644,p8645);
FA fa3470(ip_40_58,ip_41_57,ip_42_56,p8646,p8647);
FA fa3471(ip_43_55,ip_44_54,ip_45_53,p8648,p8649);
FA fa3472(ip_46_52,ip_47_51,ip_48_50,p8650,p8651);
FA fa3473(ip_49_49,ip_50_48,ip_51_47,p8652,p8653);
HA ha853(ip_52_46,ip_53_45,p8654,p8655);
FA fa3474(ip_54_44,ip_55_43,ip_56_42,p8656,p8657);
HA ha854(ip_57_41,ip_58_40,p8658,p8659);
FA fa3475(ip_59_39,ip_60_38,ip_61_37,p8660,p8661);
FA fa3476(ip_62_36,ip_63_35,p8564,p8662,p8663);
FA fa3477(p8574,p8576,p8645,p8664,p8665);
FA fa3478(p8655,p8659,p8643,p8666,p8667);
HA ha855(p8647,p8649,p8668,p8669);
FA fa3479(p8651,p8653,p8657,p8670,p8671);
FA fa3480(p8661,p8663,p8566,p8672,p8673);
HA ha856(p8568,p8570,p8674,p8675);
FA fa3481(p8572,p8578,p8580,p8676,p8677);
HA ha857(p8582,p8584,p8678,p8679);
FA fa3482(p8665,p8667,p8669,p8680,p8681);
FA fa3483(p8586,p8588,p8596,p8682,p8683);
FA fa3484(p8671,p8673,p8675,p8684,p8685);
FA fa3485(p8679,p8590,p8592,p8686,p8687);
FA fa3486(p8594,p8604,p8677,p8688,p8689);
FA fa3487(p8681,p8598,p8600,p8690,p8691);
FA fa3488(p8602,p8683,p8685,p8692,p8693);
FA fa3489(p8687,p8689,p8606,p8694,p8695);
FA fa3490(p8608,p8610,p8691,p8696,p8697);
FA fa3491(p8693,p8612,p8616,p8698,p8699);
FA fa3492(p8695,p8614,p8697,p8700,p8701);
HA ha858(p8618,p8699,p8702,p8703);
FA fa3493(p8620,p8624,p8701,p8704,p8705);
FA fa3494(p8703,p8622,p8626,p8706,p8707);
FA fa3495(p8628,p8630,p8705,p8708,p8709);
HA ha859(p8632,p8707,p8710,p8711);
FA fa3496(p8634,p8709,p8711,p8712,p8713);
FA fa3497(p8636,p8713,p8638,p8714,p8715);
HA ha860(ip_36_63,ip_37_62,p8716,p8717);
FA fa3498(ip_38_61,ip_39_60,ip_40_59,p8718,p8719);
HA ha861(ip_41_58,ip_42_57,p8720,p8721);
HA ha862(ip_43_56,ip_44_55,p8722,p8723);
FA fa3499(ip_45_54,ip_46_53,ip_47_52,p8724,p8725);
FA fa3500(ip_48_51,ip_49_50,ip_50_49,p8726,p8727);
HA ha863(ip_51_48,ip_52_47,p8728,p8729);
FA fa3501(ip_53_46,ip_54_45,ip_55_44,p8730,p8731);
FA fa3502(ip_56_43,ip_57_42,ip_58_41,p8732,p8733);
FA fa3503(ip_59_40,ip_60_39,ip_61_38,p8734,p8735);
FA fa3504(ip_62_37,ip_63_36,p8644,p8736,p8737);
FA fa3505(p8654,p8658,p8717,p8738,p8739);
FA fa3506(p8721,p8723,p8729,p8740,p8741);
HA ha864(p8719,p8725,p8742,p8743);
FA fa3507(p8727,p8731,p8733,p8744,p8745);
FA fa3508(p8735,p8737,p8642,p8746,p8747);
FA fa3509(p8646,p8648,p8650,p8748,p8749);
FA fa3510(p8652,p8656,p8660,p8750,p8751);
FA fa3511(p8662,p8668,p8739,p8752,p8753);
FA fa3512(p8741,p8743,p8664,p8754,p8755);
FA fa3513(p8666,p8674,p8678,p8756,p8757);
HA ha865(p8745,p8747,p8758,p8759);
FA fa3514(p8670,p8672,p8749,p8760,p8761);
FA fa3515(p8751,p8753,p8755,p8762,p8763);
FA fa3516(p8759,p8676,p8680,p8764,p8765);
FA fa3517(p8757,p8682,p8684,p8766,p8767);
FA fa3518(p8761,p8763,p8686,p8768,p8769);
FA fa3519(p8688,p8765,p8690,p8770,p8771);
FA fa3520(p8692,p8767,p8769,p8772,p8773);
FA fa3521(p8694,p8771,p8696,p8774,p8775);
FA fa3522(p8773,p8698,p8702,p8776,p8777);
HA ha866(p8775,p8700,p8778,p8779);
FA fa3523(p8777,p8779,p8704,p8780,p8781);
FA fa3524(p8706,p8710,p8781,p8782,p8783);
FA fa3525(p8708,p8783,p8712,p8784,p8785);
FA fa3526(ip_37_63,ip_38_62,ip_39_61,p8786,p8787);
FA fa3527(ip_40_60,ip_41_59,ip_42_58,p8788,p8789);
FA fa3528(ip_43_57,ip_44_56,ip_45_55,p8790,p8791);
FA fa3529(ip_46_54,ip_47_53,ip_48_52,p8792,p8793);
FA fa3530(ip_49_51,ip_50_50,ip_51_49,p8794,p8795);
FA fa3531(ip_52_48,ip_53_47,ip_54_46,p8796,p8797);
FA fa3532(ip_55_45,ip_56_44,ip_57_43,p8798,p8799);
FA fa3533(ip_58_42,ip_59_41,ip_60_40,p8800,p8801);
FA fa3534(ip_61_39,ip_62_38,ip_63_37,p8802,p8803);
FA fa3535(p8716,p8720,p8722,p8804,p8805);
HA ha867(p8728,p8787,p8806,p8807);
HA ha868(p8789,p8791,p8808,p8809);
HA ha869(p8793,p8795,p8810,p8811);
HA ha870(p8797,p8799,p8812,p8813);
FA fa3536(p8801,p8803,p8718,p8814,p8815);
FA fa3537(p8724,p8726,p8730,p8816,p8817);
FA fa3538(p8732,p8734,p8736,p8818,p8819);
FA fa3539(p8742,p8805,p8807,p8820,p8821);
FA fa3540(p8809,p8811,p8813,p8822,p8823);
FA fa3541(p8738,p8740,p8815,p8824,p8825);
FA fa3542(p8744,p8746,p8758,p8826,p8827);
FA fa3543(p8817,p8819,p8821,p8828,p8829);
FA fa3544(p8823,p8748,p8750,p8830,p8831);
FA fa3545(p8752,p8754,p8825,p8832,p8833);
FA fa3546(p8756,p8827,p8829,p8834,p8835);
FA fa3547(p8760,p8762,p8831,p8836,p8837);
FA fa3548(p8833,p8764,p8835,p8838,p8839);
HA ha871(p8766,p8768,p8840,p8841);
HA ha872(p8837,p8770,p8842,p8843);
FA fa3549(p8839,p8841,p8772,p8844,p8845);
FA fa3550(p8843,p8774,p8845,p8846,p8847);
FA fa3551(p8778,p8776,p8847,p8848,p8849);
FA fa3552(p8780,p8849,p8782,p8850,p8851);
HA ha873(ip_38_63,ip_39_62,p8852,p8853);
FA fa3553(ip_40_61,ip_41_60,ip_42_59,p8854,p8855);
FA fa3554(ip_43_58,ip_44_57,ip_45_56,p8856,p8857);
FA fa3555(ip_46_55,ip_47_54,ip_48_53,p8858,p8859);
FA fa3556(ip_49_52,ip_50_51,ip_51_50,p8860,p8861);
FA fa3557(ip_52_49,ip_53_48,ip_54_47,p8862,p8863);
FA fa3558(ip_55_46,ip_56_45,ip_57_44,p8864,p8865);
FA fa3559(ip_58_43,ip_59_42,ip_60_41,p8866,p8867);
FA fa3560(ip_61_40,ip_62_39,ip_63_38,p8868,p8869);
HA ha874(p8853,p8855,p8870,p8871);
FA fa3561(p8857,p8859,p8861,p8872,p8873);
FA fa3562(p8863,p8865,p8867,p8874,p8875);
FA fa3563(p8869,p8786,p8788,p8876,p8877);
FA fa3564(p8790,p8792,p8794,p8878,p8879);
FA fa3565(p8796,p8798,p8800,p8880,p8881);
FA fa3566(p8802,p8806,p8808,p8882,p8883);
FA fa3567(p8810,p8812,p8871,p8884,p8885);
HA ha875(p8804,p8873,p8886,p8887);
FA fa3568(p8875,p8814,p8877,p8888,p8889);
FA fa3569(p8879,p8881,p8883,p8890,p8891);
FA fa3570(p8885,p8887,p8816,p8892,p8893);
FA fa3571(p8818,p8820,p8822,p8894,p8895);
FA fa3572(p8824,p8889,p8891,p8896,p8897);
FA fa3573(p8893,p8826,p8828,p8898,p8899);
FA fa3574(p8895,p8830,p8832,p8900,p8901);
FA fa3575(p8897,p8834,p8899,p8902,p8903);
FA fa3576(p8836,p8840,p8901,p8904,p8905);
HA ha876(p8838,p8842,p8906,p8907);
FA fa3577(p8903,p8905,p8907,p8908,p8909);
FA fa3578(p8844,p8909,p8846,p8910,p8911);
FA fa3579(p8911,p8848,p8850,p8912,p8913);
FA fa3580(ip_39_63,ip_40_62,ip_41_61,p8914,p8915);
FA fa3581(ip_42_60,ip_43_59,ip_44_58,p8916,p8917);
FA fa3582(ip_45_57,ip_46_56,ip_47_55,p8918,p8919);
FA fa3583(ip_48_54,ip_49_53,ip_50_52,p8920,p8921);
FA fa3584(ip_51_51,ip_52_50,ip_53_49,p8922,p8923);
FA fa3585(ip_54_48,ip_55_47,ip_56_46,p8924,p8925);
FA fa3586(ip_57_45,ip_58_44,ip_59_43,p8926,p8927);
FA fa3587(ip_60_42,ip_61_41,ip_62_40,p8928,p8929);
HA ha877(ip_63_39,p8852,p8930,p8931);
HA ha878(p8915,p8917,p8932,p8933);
FA fa3588(p8919,p8921,p8923,p8934,p8935);
HA ha879(p8925,p8927,p8936,p8937);
FA fa3589(p8929,p8931,p8854,p8938,p8939);
FA fa3590(p8856,p8858,p8860,p8940,p8941);
FA fa3591(p8862,p8864,p8866,p8942,p8943);
FA fa3592(p8868,p8870,p8933,p8944,p8945);
FA fa3593(p8937,p8935,p8939,p8946,p8947);
HA ha880(p8872,p8874,p8948,p8949);
HA ha881(p8886,p8941,p8950,p8951);
FA fa3594(p8943,p8945,p8876,p8952,p8953);
FA fa3595(p8878,p8880,p8882,p8954,p8955);
FA fa3596(p8884,p8947,p8949,p8956,p8957);
FA fa3597(p8951,p8953,p8888,p8958,p8959);
FA fa3598(p8890,p8892,p8955,p8960,p8961);
FA fa3599(p8957,p8894,p8959,p8962,p8963);
FA fa3600(p8896,p8961,p8898,p8964,p8965);
HA ha882(p8963,p8900,p8966,p8967);
HA ha883(p8965,p8902,p8968,p8969);
FA fa3601(p8906,p8967,p8904,p8970,p8971);
HA ha884(p8969,p8971,p8972,p8973);
FA fa3602(p8908,p8973,p8910,p8974,p8975);
FA fa3603(ip_40_63,ip_41_62,ip_42_61,p8976,p8977);
FA fa3604(ip_43_60,ip_44_59,ip_45_58,p8978,p8979);
FA fa3605(ip_46_57,ip_47_56,ip_48_55,p8980,p8981);
FA fa3606(ip_49_54,ip_50_53,ip_51_52,p8982,p8983);
HA ha885(ip_52_51,ip_53_50,p8984,p8985);
FA fa3607(ip_54_49,ip_55_48,ip_56_47,p8986,p8987);
FA fa3608(ip_57_46,ip_58_45,ip_59_44,p8988,p8989);
FA fa3609(ip_60_43,ip_61_42,ip_62_41,p8990,p8991);
FA fa3610(ip_63_40,p8985,p8930,p8992,p8993);
FA fa3611(p8977,p8979,p8981,p8994,p8995);
FA fa3612(p8983,p8987,p8989,p8996,p8997);
FA fa3613(p8991,p8914,p8916,p8998,p8999);
FA fa3614(p8918,p8920,p8922,p9000,p9001);
FA fa3615(p8924,p8926,p8928,p9002,p9003);
HA ha886(p8932,p8936,p9004,p9005);
FA fa3616(p8993,p8995,p8997,p9006,p9007);
FA fa3617(p9005,p8934,p8938,p9008,p9009);
FA fa3618(p8999,p9001,p9003,p9010,p9011);
FA fa3619(p8940,p8942,p8944,p9012,p9013);
FA fa3620(p8948,p8950,p9007,p9014,p9015);
FA fa3621(p8946,p9009,p9011,p9016,p9017);
FA fa3622(p8952,p9013,p9015,p9018,p9019);
FA fa3623(p8954,p8956,p9017,p9020,p9021);
FA fa3624(p8958,p9019,p8960,p9022,p9023);
FA fa3625(p9021,p8962,p9023,p9024,p9025);
FA fa3626(p8964,p8966,p8968,p9026,p9027);
HA ha887(p9025,p9027,p9028,p9029);
FA fa3627(p8970,p8972,p9029,p9030,p9031);
FA fa3628(ip_41_63,ip_42_62,ip_43_61,p9032,p9033);
FA fa3629(ip_44_60,ip_45_59,ip_46_58,p9034,p9035);
HA ha888(ip_47_57,ip_48_56,p9036,p9037);
FA fa3630(ip_49_55,ip_50_54,ip_51_53,p9038,p9039);
FA fa3631(ip_52_52,ip_53_51,ip_54_50,p9040,p9041);
FA fa3632(ip_55_49,ip_56_48,ip_57_47,p9042,p9043);
FA fa3633(ip_58_46,ip_59_45,ip_60_44,p9044,p9045);
FA fa3634(ip_61_43,ip_62_42,ip_63_41,p9046,p9047);
FA fa3635(p8984,p9037,p9033,p9048,p9049);
FA fa3636(p9035,p9039,p9041,p9050,p9051);
FA fa3637(p9043,p9045,p9047,p9052,p9053);
FA fa3638(p8976,p8978,p8980,p9054,p9055);
FA fa3639(p8982,p8986,p8988,p9056,p9057);
FA fa3640(p8990,p9049,p8992,p9058,p9059);
FA fa3641(p9004,p9051,p9053,p9060,p9061);
FA fa3642(p8994,p8996,p9055,p9062,p9063);
FA fa3643(p9057,p9059,p8998,p9064,p9065);
FA fa3644(p9000,p9002,p9061,p9066,p9067);
FA fa3645(p9006,p9063,p9065,p9068,p9069);
FA fa3646(p9008,p9010,p9067,p9070,p9071);
FA fa3647(p9012,p9014,p9069,p9072,p9073);
FA fa3648(p9016,p9071,p9018,p9074,p9075);
FA fa3649(p9073,p9020,p9075,p9076,p9077);
FA fa3650(p9022,p9077,p9024,p9078,p9079);
FA fa3651(p9026,p9028,p9079,p9080,p9081);
FA fa3652(ip_42_63,ip_43_62,ip_44_61,p9082,p9083);
FA fa3653(ip_45_60,ip_46_59,ip_47_58,p9084,p9085);
FA fa3654(ip_48_57,ip_49_56,ip_50_55,p9086,p9087);
FA fa3655(ip_51_54,ip_52_53,ip_53_52,p9088,p9089);
HA ha889(ip_54_51,ip_55_50,p9090,p9091);
HA ha890(ip_56_49,ip_57_48,p9092,p9093);
HA ha891(ip_58_47,ip_59_46,p9094,p9095);
FA fa3656(ip_60_45,ip_61_44,ip_62_43,p9096,p9097);
FA fa3657(ip_63_42,p9036,p9091,p9098,p9099);
FA fa3658(p9093,p9095,p9083,p9100,p9101);
FA fa3659(p9085,p9087,p9089,p9102,p9103);
FA fa3660(p9097,p9032,p9034,p9104,p9105);
FA fa3661(p9038,p9040,p9042,p9106,p9107);
FA fa3662(p9044,p9046,p9099,p9108,p9109);
FA fa3663(p9101,p9048,p9103,p9110,p9111);
FA fa3664(p9050,p9052,p9105,p9112,p9113);
HA ha892(p9107,p9109,p9114,p9115);
FA fa3665(p9054,p9056,p9058,p9116,p9117);
FA fa3666(p9111,p9115,p9060,p9118,p9119);
HA ha893(p9113,p9062,p9120,p9121);
FA fa3667(p9064,p9117,p9119,p9122,p9123);
FA fa3668(p9066,p9121,p9068,p9124,p9125);
FA fa3669(p9123,p9070,p9125,p9126,p9127);
FA fa3670(p9072,p9074,p9127,p9128,p9129);
FA fa3671(p9076,p9129,p9078,p9130,p9131);
FA fa3672(ip_43_63,ip_44_62,ip_45_61,p9132,p9133);
HA ha894(ip_46_60,ip_47_59,p9134,p9135);
HA ha895(ip_48_58,ip_49_57,p9136,p9137);
FA fa3673(ip_50_56,ip_51_55,ip_52_54,p9138,p9139);
FA fa3674(ip_53_53,ip_54_52,ip_55_51,p9140,p9141);
FA fa3675(ip_56_50,ip_57_49,ip_58_48,p9142,p9143);
FA fa3676(ip_59_47,ip_60_46,ip_61_45,p9144,p9145);
HA ha896(ip_62_44,ip_63_43,p9146,p9147);
HA ha897(p9090,p9092,p9148,p9149);
FA fa3677(p9094,p9135,p9137,p9150,p9151);
FA fa3678(p9147,p9133,p9139,p9152,p9153);
FA fa3679(p9141,p9143,p9145,p9154,p9155);
FA fa3680(p9149,p9082,p9084,p9156,p9157);
FA fa3681(p9086,p9088,p9096,p9158,p9159);
FA fa3682(p9151,p9098,p9100,p9160,p9161);
FA fa3683(p9153,p9155,p9102,p9162,p9163);
FA fa3684(p9157,p9159,p9104,p9164,p9165);
FA fa3685(p9106,p9108,p9114,p9166,p9167);
HA ha898(p9161,p9163,p9168,p9169);
FA fa3686(p9110,p9165,p9169,p9170,p9171);
FA fa3687(p9112,p9167,p9116,p9172,p9173);
FA fa3688(p9118,p9120,p9171,p9174,p9175);
FA fa3689(p9173,p9122,p9175,p9176,p9177);
HA ha899(p9124,p9177,p9178,p9179);
HA ha900(p9126,p9179,p9180,p9181);
FA fa3690(p9181,p9128,p9130,p9182,p9183);
HA ha901(ip_44_63,ip_45_62,p9184,p9185);
HA ha902(ip_46_61,ip_47_60,p9186,p9187);
FA fa3691(ip_48_59,ip_49_58,ip_50_57,p9188,p9189);
HA ha903(ip_51_56,ip_52_55,p9190,p9191);
FA fa3692(ip_53_54,ip_54_53,ip_55_52,p9192,p9193);
FA fa3693(ip_56_51,ip_57_50,ip_58_49,p9194,p9195);
FA fa3694(ip_59_48,ip_60_47,ip_61_46,p9196,p9197);
FA fa3695(ip_62_45,ip_63_44,p9134,p9198,p9199);
FA fa3696(p9136,p9146,p9185,p9200,p9201);
FA fa3697(p9187,p9191,p9148,p9202,p9203);
HA ha904(p9189,p9193,p9204,p9205);
FA fa3698(p9195,p9197,p9199,p9206,p9207);
FA fa3699(p9132,p9138,p9140,p9208,p9209);
FA fa3700(p9142,p9144,p9201,p9210,p9211);
FA fa3701(p9203,p9205,p9150,p9212,p9213);
HA ha905(p9207,p9152,p9214,p9215);
FA fa3702(p9154,p9209,p9211,p9216,p9217);
FA fa3703(p9213,p9156,p9158,p9218,p9219);
FA fa3704(p9215,p9160,p9162,p9220,p9221);
FA fa3705(p9168,p9217,p9164,p9222,p9223);
HA ha906(p9219,p9166,p9224,p9225);
FA fa3706(p9221,p9223,p9170,p9226,p9227);
FA fa3707(p9225,p9172,p9227,p9228,p9229);
FA fa3708(p9174,p9229,p9176,p9230,p9231);
FA fa3709(p9178,p9180,p9231,p9232,p9233);
FA fa3710(ip_45_63,ip_46_62,ip_47_61,p9234,p9235);
HA ha907(ip_48_60,ip_49_59,p9236,p9237);
FA fa3711(ip_50_58,ip_51_57,ip_52_56,p9238,p9239);
HA ha908(ip_53_55,ip_54_54,p9240,p9241);
HA ha909(ip_55_53,ip_56_52,p9242,p9243);
HA ha910(ip_57_51,ip_58_50,p9244,p9245);
FA fa3712(ip_59_49,ip_60_48,ip_61_47,p9246,p9247);
HA ha911(ip_62_46,ip_63_45,p9248,p9249);
FA fa3713(p9184,p9186,p9190,p9250,p9251);
FA fa3714(p9237,p9241,p9243,p9252,p9253);
FA fa3715(p9245,p9249,p9235,p9254,p9255);
FA fa3716(p9239,p9247,p9188,p9256,p9257);
FA fa3717(p9192,p9194,p9196,p9258,p9259);
FA fa3718(p9198,p9204,p9251,p9260,p9261);
FA fa3719(p9253,p9255,p9200,p9262,p9263);
FA fa3720(p9202,p9257,p9206,p9264,p9265);
HA ha912(p9259,p9261,p9266,p9267);
FA fa3721(p9263,p9208,p9210,p9268,p9269);
HA ha913(p9212,p9214,p9270,p9271);
FA fa3722(p9265,p9267,p9271,p9272,p9273);
FA fa3723(p9216,p9269,p9273,p9274,p9275);
FA fa3724(p9218,p9220,p9222,p9276,p9277);
HA ha914(p9224,p9275,p9278,p9279);
HA ha915(p9279,p9226,p9280,p9281);
FA fa3725(p9277,p9281,p9228,p9282,p9283);
HA ha916(p9283,p9230,p9284,p9285);
FA fa3726(ip_46_63,ip_47_62,ip_48_61,p9286,p9287);
FA fa3727(ip_49_60,ip_50_59,ip_51_58,p9288,p9289);
FA fa3728(ip_52_57,ip_53_56,ip_54_55,p9290,p9291);
FA fa3729(ip_55_54,ip_56_53,ip_57_52,p9292,p9293);
FA fa3730(ip_58_51,ip_59_50,ip_60_49,p9294,p9295);
FA fa3731(ip_61_48,ip_62_47,ip_63_46,p9296,p9297);
FA fa3732(p9236,p9240,p9242,p9298,p9299);
HA ha917(p9244,p9248,p9300,p9301);
FA fa3733(p9287,p9289,p9291,p9302,p9303);
FA fa3734(p9293,p9295,p9297,p9304,p9305);
FA fa3735(p9301,p9234,p9238,p9306,p9307);
HA ha918(p9246,p9299,p9308,p9309);
FA fa3736(p9250,p9252,p9254,p9310,p9311);
FA fa3737(p9303,p9305,p9309,p9312,p9313);
FA fa3738(p9256,p9307,p9258,p9314,p9315);
FA fa3739(p9260,p9262,p9266,p9316,p9317);
HA ha919(p9311,p9313,p9318,p9319);
HA ha920(p9264,p9270,p9320,p9321);
FA fa3740(p9315,p9319,p9317,p9322,p9323);
HA ha921(p9321,p9268,p9324,p9325);
FA fa3741(p9272,p9323,p9325,p9326,p9327);
FA fa3742(p9274,p9278,p9327,p9328,p9329);
FA fa3743(p9276,p9280,p9329,p9330,p9331);
FA fa3744(p9331,p9282,p9284,p9332,p9333);
FA fa3745(ip_47_63,ip_48_62,ip_49_61,p9334,p9335);
HA ha922(ip_50_60,ip_51_59,p9336,p9337);
HA ha923(ip_52_58,ip_53_57,p9338,p9339);
FA fa3746(ip_54_56,ip_55_55,ip_56_54,p9340,p9341);
HA ha924(ip_57_53,ip_58_52,p9342,p9343);
HA ha925(ip_59_51,ip_60_50,p9344,p9345);
FA fa3747(ip_61_49,ip_62_48,ip_63_47,p9346,p9347);
FA fa3748(p9337,p9339,p9343,p9348,p9349);
FA fa3749(p9345,p9300,p9335,p9350,p9351);
FA fa3750(p9341,p9347,p9286,p9352,p9353);
FA fa3751(p9288,p9290,p9292,p9354,p9355);
FA fa3752(p9294,p9296,p9349,p9356,p9357);
FA fa3753(p9298,p9308,p9351,p9358,p9359);
FA fa3754(p9353,p9302,p9304,p9360,p9361);
FA fa3755(p9355,p9357,p9306,p9362,p9363);
FA fa3756(p9359,p9310,p9312,p9364,p9365);
FA fa3757(p9318,p9361,p9363,p9366,p9367);
FA fa3758(p9314,p9320,p9316,p9368,p9369);
HA ha926(p9365,p9367,p9370,p9371);
FA fa3759(p9322,p9324,p9369,p9372,p9373);
FA fa3760(p9371,p9326,p9373,p9374,p9375);
FA fa3761(p9328,p9375,p9330,p9376,p9377);
FA fa3762(ip_48_63,ip_49_62,ip_50_61,p9378,p9379);
FA fa3763(ip_51_60,ip_52_59,ip_53_58,p9380,p9381);
FA fa3764(ip_54_57,ip_55_56,ip_56_55,p9382,p9383);
HA ha927(ip_57_54,ip_58_53,p9384,p9385);
FA fa3765(ip_59_52,ip_60_51,ip_61_50,p9386,p9387);
HA ha928(ip_62_49,ip_63_48,p9388,p9389);
FA fa3766(p9336,p9338,p9342,p9390,p9391);
FA fa3767(p9344,p9385,p9389,p9392,p9393);
FA fa3768(p9379,p9381,p9383,p9394,p9395);
FA fa3769(p9387,p9334,p9340,p9396,p9397);
HA ha929(p9346,p9391,p9398,p9399);
HA ha930(p9393,p9348,p9400,p9401);
FA fa3770(p9395,p9399,p9350,p9402,p9403);
FA fa3771(p9352,p9397,p9401,p9404,p9405);
FA fa3772(p9354,p9356,p9403,p9406,p9407);
FA fa3773(p9358,p9405,p9360,p9408,p9409);
FA fa3774(p9362,p9407,p9409,p9410,p9411);
FA fa3775(p9364,p9366,p9370,p9412,p9413);
HA ha931(p9411,p9368,p9414,p9415);
FA fa3776(p9413,p9415,p9372,p9416,p9417);
FA fa3777(p9417,p9374,p9376,p9418,p9419);
FA fa3778(ip_49_63,ip_50_62,ip_51_61,p9420,p9421);
FA fa3779(ip_52_60,ip_53_59,ip_54_58,p9422,p9423);
FA fa3780(ip_55_57,ip_56_56,ip_57_55,p9424,p9425);
HA ha932(ip_58_54,ip_59_53,p9426,p9427);
HA ha933(ip_60_52,ip_61_51,p9428,p9429);
FA fa3781(ip_62_50,ip_63_49,p9384,p9430,p9431);
FA fa3782(p9388,p9427,p9429,p9432,p9433);
FA fa3783(p9421,p9423,p9425,p9434,p9435);
FA fa3784(p9431,p9378,p9380,p9436,p9437);
FA fa3785(p9382,p9386,p9433,p9438,p9439);
FA fa3786(p9390,p9392,p9398,p9440,p9441);
FA fa3787(p9435,p9394,p9400,p9442,p9443);
HA ha934(p9437,p9439,p9444,p9445);
FA fa3788(p9396,p9441,p9445,p9446,p9447);
FA fa3789(p9402,p9443,p9404,p9448,p9449);
FA fa3790(p9447,p9406,p9449,p9450,p9451);
HA ha935(p9408,p9410,p9452,p9453);
FA fa3791(p9451,p9414,p9453,p9454,p9455);
FA fa3792(p9412,p9455,p9416,p9456,p9457);
FA fa3793(ip_50_63,ip_51_62,ip_52_61,p9458,p9459);
FA fa3794(ip_53_60,ip_54_59,ip_55_58,p9460,p9461);
HA ha936(ip_56_57,ip_57_56,p9462,p9463);
FA fa3795(ip_58_55,ip_59_54,ip_60_53,p9464,p9465);
FA fa3796(ip_61_52,ip_62_51,ip_63_50,p9466,p9467);
FA fa3797(p9426,p9428,p9463,p9468,p9469);
FA fa3798(p9459,p9461,p9465,p9470,p9471);
HA ha937(p9467,p9420,p9472,p9473);
FA fa3799(p9422,p9424,p9430,p9474,p9475);
FA fa3800(p9469,p9432,p9471,p9476,p9477);
FA fa3801(p9473,p9434,p9475,p9478,p9479);
FA fa3802(p9436,p9438,p9444,p9480,p9481);
FA fa3803(p9477,p9440,p9479,p9482,p9483);
FA fa3804(p9442,p9481,p9446,p9484,p9485);
FA fa3805(p9483,p9448,p9485,p9486,p9487);
FA fa3806(p9450,p9452,p9487,p9488,p9489);
FA fa3807(p9489,p9454,p9456,p9490,p9491);
FA fa3808(ip_51_63,ip_52_62,ip_53_61,p9492,p9493);
HA ha938(ip_54_60,ip_55_59,p9494,p9495);
FA fa3809(ip_56_58,ip_57_57,ip_58_56,p9496,p9497);
FA fa3810(ip_59_55,ip_60_54,ip_61_53,p9498,p9499);
FA fa3811(ip_62_52,ip_63_51,p9462,p9500,p9501);
HA ha939(p9495,p9493,p9502,p9503);
FA fa3812(p9497,p9499,p9501,p9504,p9505);
FA fa3813(p9458,p9460,p9464,p9506,p9507);
FA fa3814(p9466,p9503,p9468,p9508,p9509);
FA fa3815(p9472,p9505,p9470,p9510,p9511);
FA fa3816(p9507,p9509,p9474,p9512,p9513);
FA fa3817(p9511,p9476,p9513,p9514,p9515);
FA fa3818(p9478,p9480,p9515,p9516,p9517);
FA fa3819(p9482,p9484,p9517,p9518,p9519);
FA fa3820(p9486,p9519,p9488,p9520,p9521);
FA fa3821(ip_52_63,ip_53_62,ip_54_61,p9522,p9523);
FA fa3822(ip_55_60,ip_56_59,ip_57_58,p9524,p9525);
HA ha940(ip_58_57,ip_59_56,p9526,p9527);
FA fa3823(ip_60_55,ip_61_54,ip_62_53,p9528,p9529);
FA fa3824(ip_63_52,p9494,p9527,p9530,p9531);
FA fa3825(p9523,p9525,p9529,p9532,p9533);
FA fa3826(p9492,p9496,p9498,p9534,p9535);
HA ha941(p9500,p9502,p9536,p9537);
FA fa3827(p9531,p9533,p9537,p9538,p9539);
FA fa3828(p9504,p9535,p9506,p9540,p9541);
HA ha942(p9508,p9539,p9542,p9543);
FA fa3829(p9510,p9541,p9543,p9544,p9545);
FA fa3830(p9512,p9545,p9514,p9546,p9547);
FA fa3831(p9547,p9516,p9518,p9548,p9549);
FA fa3832(ip_53_63,ip_54_62,ip_55_61,p9550,p9551);
FA fa3833(ip_56_60,ip_57_59,ip_58_58,p9552,p9553);
FA fa3834(ip_59_57,ip_60_56,ip_61_55,p9554,p9555);
HA ha943(ip_62_54,ip_63_53,p9556,p9557);
HA ha944(p9526,p9557,p9558,p9559);
FA fa3835(p9551,p9553,p9555,p9560,p9561);
FA fa3836(p9559,p9522,p9524,p9562,p9563);
FA fa3837(p9528,p9530,p9536,p9564,p9565);
HA ha945(p9561,p9532,p9566,p9567);
HA ha946(p9563,p9534,p9568,p9569);
HA ha947(p9565,p9567,p9570,p9571);
HA ha948(p9538,p9542,p9572,p9573);
FA fa3838(p9569,p9571,p9540,p9574,p9575);
FA fa3839(p9573,p9575,p9544,p9576,p9577);
FA fa3840(p9577,p9546,p9548,p9578,p9579);
FA fa3841(ip_54_63,ip_55_62,ip_56_61,p9580,p9581);
FA fa3842(ip_57_60,ip_58_59,ip_59_58,p9582,p9583);
FA fa3843(ip_60_57,ip_61_56,ip_62_55,p9584,p9585);
FA fa3844(ip_63_54,p9556,p9558,p9586,p9587);
FA fa3845(p9581,p9583,p9585,p9588,p9589);
FA fa3846(p9550,p9552,p9554,p9590,p9591);
FA fa3847(p9587,p9589,p9560,p9592,p9593);
FA fa3848(p9591,p9562,p9566,p9594,p9595);
FA fa3849(p9593,p9564,p9568,p9596,p9597);
FA fa3850(p9570,p9572,p9595,p9598,p9599);
FA fa3851(p9597,p9574,p9599,p9600,p9601);
FA fa3852(p9576,p9601,p9578,p9602,p9603);
FA fa3853(ip_55_63,ip_56_62,ip_57_61,p9604,p9605);
HA ha949(ip_58_60,ip_59_59,p9606,p9607);
FA fa3854(ip_60_58,ip_61_57,ip_62_56,p9608,p9609);
FA fa3855(ip_63_55,p9607,p9605,p9610,p9611);
FA fa3856(p9609,p9580,p9582,p9612,p9613);
FA fa3857(p9584,p9611,p9586,p9614,p9615);
FA fa3858(p9588,p9613,p9615,p9616,p9617);
FA fa3859(p9590,p9592,p9617,p9618,p9619);
HA ha950(p9594,p9619,p9620,p9621);
FA fa3860(p9596,p9621,p9598,p9622,p9623);
FA fa3861(p9623,p9600,p9602,p9624,p9625);
FA fa3862(ip_56_63,ip_57_62,ip_58_61,p9626,p9627);
FA fa3863(ip_59_60,ip_60_59,ip_61_58,p9628,p9629);
FA fa3864(ip_62_57,ip_63_56,p9606,p9630,p9631);
FA fa3865(p9627,p9629,p9631,p9632,p9633);
FA fa3866(p9604,p9608,p9610,p9634,p9635);
FA fa3867(p9633,p9635,p9612,p9636,p9637);
FA fa3868(p9614,p9637,p9616,p9638,p9639);
FA fa3869(p9639,p9618,p9620,p9640,p9641);
FA fa3870(p9641,p9622,p9624,p9642,p9643);
FA fa3871(ip_57_63,ip_58_62,ip_59_61,p9644,p9645);
FA fa3872(ip_60_60,ip_61_59,ip_62_58,p9646,p9647);
FA fa3873(ip_63_57,p9645,p9647,p9648,p9649);
FA fa3874(p9626,p9628,p9630,p9650,p9651);
HA ha951(p9649,p9632,p9652,p9653);
FA fa3875(p9651,p9634,p9653,p9654,p9655);
FA fa3876(p9636,p9655,p9638,p9656,p9657);
FA fa3877(p9657,p9640,p9642,p9658,p9659);
FA fa3878(ip_58_63,ip_59_62,ip_60_61,p9660,p9661);
FA fa3879(ip_61_60,ip_62_59,ip_63_58,p9662,p9663);
FA fa3880(p9661,p9663,p9644,p9664,p9665);
FA fa3881(p9646,p9665,p9648,p9666,p9667);
FA fa3882(p9650,p9652,p9667,p9668,p9669);
FA fa3883(p9669,p9654,p9656,p9670,p9671);
FA fa3884(ip_59_63,ip_60_62,ip_61_61,p9672,p9673);
HA ha952(ip_62_60,ip_63_59,p9674,p9675);
FA fa3885(p9675,p9673,p9660,p9676,p9677);
HA ha953(p9662,p9677,p9678,p9679);
FA fa3886(p9664,p9679,p9666,p9680,p9681);
FA fa3887(p9681,p9668,p9670,p9682,p9683);
FA fa3888(ip_60_63,ip_61_62,ip_62_61,p9684,p9685);
FA fa3889(ip_63_60,p9674,p9685,p9686,p9687);
HA ha954(p9672,p9687,p9688,p9689);
FA fa3890(p9689,p9676,p9678,p9690,p9691);
FA fa3891(p9691,p9680,p9682,p9692,p9693);
FA fa3892(ip_61_63,ip_62_62,ip_63_61,p9694,p9695);
FA fa3893(p9695,p9684,p9686,p9696,p9697);
FA fa3894(p9688,p9697,p9690,p9698,p9699);
FA fa3895(ip_62_63,ip_63_62,p9694,p9700,p9701);
FA fa3896(p9701,p9696,p9698,p9702,p9703);
HA ha955(ip_63_63,p9700,p9704,p9705);
wire [127:0] a,b;
wire [127:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = ip_2_0;
assign b[2] = p1;
assign a[3] = p3;
assign b[3] = p5;
assign a[4] = p2;
assign b[4] = p11;
assign a[5] = p10;
assign b[5] = p19;
assign a[6] = p18;
assign b[6] = p29;
assign a[7] = p28;
assign b[7] = p43;
assign a[8] = p59;
assign b[8] = 1'b0;
assign a[9] = p77;
assign b[9] = p58;
assign a[10] = p99;
assign b[10] = 1'b0;
assign a[11] = p125;
assign b[11] = 1'b0;
assign a[12] = p155;
assign b[12] = 1'b0;
assign a[13] = p185;
assign b[13] = p154;
assign a[14] = p215;
assign b[14] = 1'b0;
assign a[15] = p247;
assign b[15] = p214;
assign a[16] = p281;
assign b[16] = p246;
assign a[17] = p319;
assign b[17] = p280;
assign a[18] = p361;
assign b[18] = 1'b0;
assign a[19] = p401;
assign b[19] = p360;
assign a[20] = p447;
assign b[20] = p400;
assign a[21] = p497;
assign b[21] = 1'b0;
assign a[22] = p551;
assign b[22] = p496;
assign a[23] = p605;
assign b[23] = 1'b0;
assign a[24] = p661;
assign b[24] = p604;
assign a[25] = p717;
assign b[25] = p660;
assign a[26] = p773;
assign b[26] = p716;
assign a[27] = p835;
assign b[27] = 1'b0;
assign a[28] = p901;
assign b[28] = p834;
assign a[29] = p971;
assign b[29] = 1'b0;
assign a[30] = p1045;
assign b[30] = 1'b0;
assign a[31] = p1117;
assign b[31] = 1'b0;
assign a[32] = p1193;
assign b[32] = p1116;
assign a[33] = p1271;
assign b[33] = p1192;
assign a[34] = p1353;
assign b[34] = p1270;
assign a[35] = p1437;
assign b[35] = p1352;
assign a[36] = p1436;
assign b[36] = p1525;
assign a[37] = p1615;
assign b[37] = 1'b0;
assign a[38] = p1703;
assign b[38] = p1614;
assign a[39] = p1791;
assign b[39] = 1'b0;
assign a[40] = p1877;
assign b[40] = p1790;
assign a[41] = p1971;
assign b[41] = p1876;
assign a[42] = p2069;
assign b[42] = 1'b0;
assign a[43] = p2169;
assign b[43] = p2068;
assign a[44] = p2168;
assign b[44] = p2273;
assign a[45] = p2377;
assign b[45] = 1'b0;
assign a[46] = p2489;
assign b[46] = p2376;
assign a[47] = p2597;
assign b[47] = p2488;
assign a[48] = p2711;
assign b[48] = 1'b0;
assign a[49] = p2827;
assign b[49] = 1'b0;
assign a[50] = p2949;
assign b[50] = 1'b0;
assign a[51] = p3065;
assign b[51] = 1'b0;
assign a[52] = p3183;
assign b[52] = p3064;
assign a[53] = p3303;
assign b[53] = p3182;
assign a[54] = p3302;
assign b[54] = p3429;
assign a[55] = p3561;
assign b[55] = 1'b0;
assign a[56] = p3699;
assign b[56] = 1'b0;
assign a[57] = p3839;
assign b[57] = 1'b0;
assign a[58] = p3985;
assign b[58] = p3838;
assign a[59] = p4135;
assign b[59] = 1'b0;
assign a[60] = p4281;
assign b[60] = p4134;
assign a[61] = p4427;
assign b[61] = 1'b0;
assign a[62] = p4575;
assign b[62] = 1'b0;
assign a[63] = p4727;
assign b[63] = 1'b0;
assign a[64] = p4883;
assign b[64] = 1'b0;
assign a[65] = p5037;
assign b[65] = 1'b0;
assign a[66] = p5191;
assign b[66] = p5036;
assign a[67] = p5345;
assign b[67] = p5190;
assign a[68] = p5493;
assign b[68] = p5344;
assign a[69] = p5641;
assign b[69] = 1'b0;
assign a[70] = p5797;
assign b[70] = 1'b0;
assign a[71] = p5941;
assign b[71] = 1'b0;
assign a[72] = p6077;
assign b[72] = 1'b0;
assign a[73] = p6215;
assign b[73] = p6076;
assign a[74] = p6349;
assign b[74] = p6214;
assign a[75] = p6479;
assign b[75] = 1'b0;
assign a[76] = p6611;
assign b[76] = p6478;
assign a[77] = p6737;
assign b[77] = 1'b0;
assign a[78] = p6867;
assign b[78] = p6736;
assign a[79] = p6989;
assign b[79] = 1'b0;
assign a[80] = p7107;
assign b[80] = p6988;
assign a[81] = p7215;
assign b[81] = p7106;
assign a[82] = p7321;
assign b[82] = p7214;
assign a[83] = p7425;
assign b[83] = p7320;
assign a[84] = p7523;
assign b[84] = p7424;
assign a[85] = p7623;
assign b[85] = p7522;
assign a[86] = p7622;
assign b[86] = p7719;
assign a[87] = p7809;
assign b[87] = p7718;
assign a[88] = p7901;
assign b[88] = 1'b0;
assign a[89] = p7991;
assign b[89] = 1'b0;
assign a[90] = p8077;
assign b[90] = p7990;
assign a[91] = p8165;
assign b[91] = p8076;
assign a[92] = p8249;
assign b[92] = 1'b0;
assign a[93] = p8335;
assign b[93] = 1'b0;
assign a[94] = p8413;
assign b[94] = p8334;
assign a[95] = p8491;
assign b[95] = 1'b0;
assign a[96] = p8563;
assign b[96] = p8490;
assign a[97] = p8641;
assign b[97] = 1'b0;
assign a[98] = p8715;
assign b[98] = p8640;
assign a[99] = p8785;
assign b[99] = p8714;
assign a[100] = p8851;
assign b[100] = p8784;
assign a[101] = p8913;
assign b[101] = 1'b0;
assign a[102] = p8975;
assign b[102] = p8912;
assign a[103] = p9031;
assign b[103] = p8974;
assign a[104] = p9081;
assign b[104] = p9030;
assign a[105] = p9131;
assign b[105] = p9080;
assign a[106] = p9183;
assign b[106] = 1'b0;
assign a[107] = p9233;
assign b[107] = p9182;
assign a[108] = p9285;
assign b[108] = p9232;
assign a[109] = p9333;
assign b[109] = 1'b0;
assign a[110] = p9377;
assign b[110] = p9332;
assign a[111] = p9419;
assign b[111] = 1'b0;
assign a[112] = p9457;
assign b[112] = p9418;
assign a[113] = p9491;
assign b[113] = 1'b0;
assign a[114] = p9521;
assign b[114] = p9490;
assign a[115] = p9549;
assign b[115] = p9520;
assign a[116] = p9579;
assign b[116] = 1'b0;
assign a[117] = p9603;
assign b[117] = 1'b0;
assign a[118] = p9625;
assign b[118] = 1'b0;
assign a[119] = p9643;
assign b[119] = 1'b0;
assign a[120] = p9659;
assign b[120] = 1'b0;
assign a[121] = p9671;
assign b[121] = p9658;
assign a[122] = p9683;
assign b[122] = 1'b0;
assign a[123] = p9693;
assign b[123] = 1'b0;
assign a[124] = p9699;
assign b[124] = p9692;
assign a[125] = p9703;
assign b[125] = 1'b0;
assign a[126] = p9705;
assign b[126] = p9702;
assign a[127] = p9704;
assign b[127] = 1'b0;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[127] = s[127];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
assign o[31] = s[31];
assign o[32] = s[32];
assign o[33] = s[33];
assign o[34] = s[34];
assign o[35] = s[35];
assign o[36] = s[36];
assign o[37] = s[37];
assign o[38] = s[38];
assign o[39] = s[39];
assign o[40] = s[40];
assign o[41] = s[41];
assign o[42] = s[42];
assign o[43] = s[43];
assign o[44] = s[44];
assign o[45] = s[45];
assign o[46] = s[46];
assign o[47] = s[47];
assign o[48] = s[48];
assign o[49] = s[49];
assign o[50] = s[50];
assign o[51] = s[51];
assign o[52] = s[52];
assign o[53] = s[53];
assign o[54] = s[54];
assign o[55] = s[55];
assign o[56] = s[56];
assign o[57] = s[57];
assign o[58] = s[58];
assign o[59] = s[59];
assign o[60] = s[60];
assign o[61] = s[61];
assign o[62] = s[62];
assign o[63] = s[63];
assign o[64] = s[64];
assign o[65] = s[65];
assign o[66] = s[66];
assign o[67] = s[67];
assign o[68] = s[68];
assign o[69] = s[69];
assign o[70] = s[70];
assign o[71] = s[71];
assign o[72] = s[72];
assign o[73] = s[73];
assign o[74] = s[74];
assign o[75] = s[75];
assign o[76] = s[76];
assign o[77] = s[77];
assign o[78] = s[78];
assign o[79] = s[79];
assign o[80] = s[80];
assign o[81] = s[81];
assign o[82] = s[82];
assign o[83] = s[83];
assign o[84] = s[84];
assign o[85] = s[85];
assign o[86] = s[86];
assign o[87] = s[87];
assign o[88] = s[88];
assign o[89] = s[89];
assign o[90] = s[90];
assign o[91] = s[91];
assign o[92] = s[92];
assign o[93] = s[93];
assign o[94] = s[94];
assign o[95] = s[95];
assign o[96] = s[96];
assign o[97] = s[97];
assign o[98] = s[98];
assign o[99] = s[99];
assign o[100] = s[100];
assign o[101] = s[101];
assign o[102] = s[102];
assign o[103] = s[103];
assign o[104] = s[104];
assign o[105] = s[105];
assign o[106] = s[106];
assign o[107] = s[107];
assign o[108] = s[108];
assign o[109] = s[109];
assign o[110] = s[110];
assign o[111] = s[111];
assign o[112] = s[112];
assign o[113] = s[113];
assign o[114] = s[114];
assign o[115] = s[115];
assign o[116] = s[116];
assign o[117] = s[117];
assign o[118] = s[118];
assign o[119] = s[119];
assign o[120] = s[120];
assign o[121] = s[121];
assign o[122] = s[122];
assign o[123] = s[123];
assign o[124] = s[124];
assign o[125] = s[125];
assign o[126] = s[126];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [127:0] a,b;
output [127:0] s;
assign s = a+b;
endmodule
