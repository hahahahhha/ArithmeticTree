// 1 2 2 1 1 1 1 2 1 1 2 2 2 2 2 2 1 2 1 2 1 2 1 1 2 2 2 1 2 1 2 1 1 2 2 2 2 2 1 2 1 2 1 2 2 1 2 1 2 2 2 2 2 2 2 1 2 2 2 1 2 2 1 2 1 1 1 2 1 2 2 1 2 1 1 2 1 1 1 1 2 2 1 1 1 1 1 2 2 1 1 2 2 1 2 2 2 2 2 2 1 2 1 2 2 2 2 1 1 2 1 2 2 2 2 1 2 2 2 2 2 2 2 2 2 2 2 2 

module main(x,y,o);
input [63:0] x,y;
output [127:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_0_8,ip_0_9,ip_0_10,ip_0_11,ip_0_12,ip_0_13,ip_0_14,ip_0_15,ip_0_16,ip_0_17,ip_0_18,ip_0_19,ip_0_20,ip_0_21,ip_0_22,ip_0_23,ip_0_24,ip_0_25,ip_0_26,ip_0_27,ip_0_28,ip_0_29,ip_0_30,ip_0_31,ip_0_32,ip_0_33,ip_0_34,ip_0_35,ip_0_36,ip_0_37,ip_0_38,ip_0_39,ip_0_40,ip_0_41,ip_0_42,ip_0_43,ip_0_44,ip_0_45,ip_0_46,ip_0_47,ip_0_48,ip_0_49,ip_0_50,ip_0_51,ip_0_52,ip_0_53,ip_0_54,ip_0_55,ip_0_56,ip_0_57,ip_0_58,ip_0_59,ip_0_60,ip_0_61,ip_0_62,ip_0_63,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_1_8,ip_1_9,ip_1_10,ip_1_11,ip_1_12,ip_1_13,ip_1_14,ip_1_15,ip_1_16,ip_1_17,ip_1_18,ip_1_19,ip_1_20,ip_1_21,ip_1_22,ip_1_23,ip_1_24,ip_1_25,ip_1_26,ip_1_27,ip_1_28,ip_1_29,ip_1_30,ip_1_31,ip_1_32,ip_1_33,ip_1_34,ip_1_35,ip_1_36,ip_1_37,ip_1_38,ip_1_39,ip_1_40,ip_1_41,ip_1_42,ip_1_43,ip_1_44,ip_1_45,ip_1_46,ip_1_47,ip_1_48,ip_1_49,ip_1_50,ip_1_51,ip_1_52,ip_1_53,ip_1_54,ip_1_55,ip_1_56,ip_1_57,ip_1_58,ip_1_59,ip_1_60,ip_1_61,ip_1_62,ip_1_63,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_2_8,ip_2_9,ip_2_10,ip_2_11,ip_2_12,ip_2_13,ip_2_14,ip_2_15,ip_2_16,ip_2_17,ip_2_18,ip_2_19,ip_2_20,ip_2_21,ip_2_22,ip_2_23,ip_2_24,ip_2_25,ip_2_26,ip_2_27,ip_2_28,ip_2_29,ip_2_30,ip_2_31,ip_2_32,ip_2_33,ip_2_34,ip_2_35,ip_2_36,ip_2_37,ip_2_38,ip_2_39,ip_2_40,ip_2_41,ip_2_42,ip_2_43,ip_2_44,ip_2_45,ip_2_46,ip_2_47,ip_2_48,ip_2_49,ip_2_50,ip_2_51,ip_2_52,ip_2_53,ip_2_54,ip_2_55,ip_2_56,ip_2_57,ip_2_58,ip_2_59,ip_2_60,ip_2_61,ip_2_62,ip_2_63,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_3_8,ip_3_9,ip_3_10,ip_3_11,ip_3_12,ip_3_13,ip_3_14,ip_3_15,ip_3_16,ip_3_17,ip_3_18,ip_3_19,ip_3_20,ip_3_21,ip_3_22,ip_3_23,ip_3_24,ip_3_25,ip_3_26,ip_3_27,ip_3_28,ip_3_29,ip_3_30,ip_3_31,ip_3_32,ip_3_33,ip_3_34,ip_3_35,ip_3_36,ip_3_37,ip_3_38,ip_3_39,ip_3_40,ip_3_41,ip_3_42,ip_3_43,ip_3_44,ip_3_45,ip_3_46,ip_3_47,ip_3_48,ip_3_49,ip_3_50,ip_3_51,ip_3_52,ip_3_53,ip_3_54,ip_3_55,ip_3_56,ip_3_57,ip_3_58,ip_3_59,ip_3_60,ip_3_61,ip_3_62,ip_3_63,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_4_8,ip_4_9,ip_4_10,ip_4_11,ip_4_12,ip_4_13,ip_4_14,ip_4_15,ip_4_16,ip_4_17,ip_4_18,ip_4_19,ip_4_20,ip_4_21,ip_4_22,ip_4_23,ip_4_24,ip_4_25,ip_4_26,ip_4_27,ip_4_28,ip_4_29,ip_4_30,ip_4_31,ip_4_32,ip_4_33,ip_4_34,ip_4_35,ip_4_36,ip_4_37,ip_4_38,ip_4_39,ip_4_40,ip_4_41,ip_4_42,ip_4_43,ip_4_44,ip_4_45,ip_4_46,ip_4_47,ip_4_48,ip_4_49,ip_4_50,ip_4_51,ip_4_52,ip_4_53,ip_4_54,ip_4_55,ip_4_56,ip_4_57,ip_4_58,ip_4_59,ip_4_60,ip_4_61,ip_4_62,ip_4_63,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_5_8,ip_5_9,ip_5_10,ip_5_11,ip_5_12,ip_5_13,ip_5_14,ip_5_15,ip_5_16,ip_5_17,ip_5_18,ip_5_19,ip_5_20,ip_5_21,ip_5_22,ip_5_23,ip_5_24,ip_5_25,ip_5_26,ip_5_27,ip_5_28,ip_5_29,ip_5_30,ip_5_31,ip_5_32,ip_5_33,ip_5_34,ip_5_35,ip_5_36,ip_5_37,ip_5_38,ip_5_39,ip_5_40,ip_5_41,ip_5_42,ip_5_43,ip_5_44,ip_5_45,ip_5_46,ip_5_47,ip_5_48,ip_5_49,ip_5_50,ip_5_51,ip_5_52,ip_5_53,ip_5_54,ip_5_55,ip_5_56,ip_5_57,ip_5_58,ip_5_59,ip_5_60,ip_5_61,ip_5_62,ip_5_63,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_6_8,ip_6_9,ip_6_10,ip_6_11,ip_6_12,ip_6_13,ip_6_14,ip_6_15,ip_6_16,ip_6_17,ip_6_18,ip_6_19,ip_6_20,ip_6_21,ip_6_22,ip_6_23,ip_6_24,ip_6_25,ip_6_26,ip_6_27,ip_6_28,ip_6_29,ip_6_30,ip_6_31,ip_6_32,ip_6_33,ip_6_34,ip_6_35,ip_6_36,ip_6_37,ip_6_38,ip_6_39,ip_6_40,ip_6_41,ip_6_42,ip_6_43,ip_6_44,ip_6_45,ip_6_46,ip_6_47,ip_6_48,ip_6_49,ip_6_50,ip_6_51,ip_6_52,ip_6_53,ip_6_54,ip_6_55,ip_6_56,ip_6_57,ip_6_58,ip_6_59,ip_6_60,ip_6_61,ip_6_62,ip_6_63,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7,ip_7_8,ip_7_9,ip_7_10,ip_7_11,ip_7_12,ip_7_13,ip_7_14,ip_7_15,ip_7_16,ip_7_17,ip_7_18,ip_7_19,ip_7_20,ip_7_21,ip_7_22,ip_7_23,ip_7_24,ip_7_25,ip_7_26,ip_7_27,ip_7_28,ip_7_29,ip_7_30,ip_7_31,ip_7_32,ip_7_33,ip_7_34,ip_7_35,ip_7_36,ip_7_37,ip_7_38,ip_7_39,ip_7_40,ip_7_41,ip_7_42,ip_7_43,ip_7_44,ip_7_45,ip_7_46,ip_7_47,ip_7_48,ip_7_49,ip_7_50,ip_7_51,ip_7_52,ip_7_53,ip_7_54,ip_7_55,ip_7_56,ip_7_57,ip_7_58,ip_7_59,ip_7_60,ip_7_61,ip_7_62,ip_7_63,ip_8_0,ip_8_1,ip_8_2,ip_8_3,ip_8_4,ip_8_5,ip_8_6,ip_8_7,ip_8_8,ip_8_9,ip_8_10,ip_8_11,ip_8_12,ip_8_13,ip_8_14,ip_8_15,ip_8_16,ip_8_17,ip_8_18,ip_8_19,ip_8_20,ip_8_21,ip_8_22,ip_8_23,ip_8_24,ip_8_25,ip_8_26,ip_8_27,ip_8_28,ip_8_29,ip_8_30,ip_8_31,ip_8_32,ip_8_33,ip_8_34,ip_8_35,ip_8_36,ip_8_37,ip_8_38,ip_8_39,ip_8_40,ip_8_41,ip_8_42,ip_8_43,ip_8_44,ip_8_45,ip_8_46,ip_8_47,ip_8_48,ip_8_49,ip_8_50,ip_8_51,ip_8_52,ip_8_53,ip_8_54,ip_8_55,ip_8_56,ip_8_57,ip_8_58,ip_8_59,ip_8_60,ip_8_61,ip_8_62,ip_8_63,ip_9_0,ip_9_1,ip_9_2,ip_9_3,ip_9_4,ip_9_5,ip_9_6,ip_9_7,ip_9_8,ip_9_9,ip_9_10,ip_9_11,ip_9_12,ip_9_13,ip_9_14,ip_9_15,ip_9_16,ip_9_17,ip_9_18,ip_9_19,ip_9_20,ip_9_21,ip_9_22,ip_9_23,ip_9_24,ip_9_25,ip_9_26,ip_9_27,ip_9_28,ip_9_29,ip_9_30,ip_9_31,ip_9_32,ip_9_33,ip_9_34,ip_9_35,ip_9_36,ip_9_37,ip_9_38,ip_9_39,ip_9_40,ip_9_41,ip_9_42,ip_9_43,ip_9_44,ip_9_45,ip_9_46,ip_9_47,ip_9_48,ip_9_49,ip_9_50,ip_9_51,ip_9_52,ip_9_53,ip_9_54,ip_9_55,ip_9_56,ip_9_57,ip_9_58,ip_9_59,ip_9_60,ip_9_61,ip_9_62,ip_9_63,ip_10_0,ip_10_1,ip_10_2,ip_10_3,ip_10_4,ip_10_5,ip_10_6,ip_10_7,ip_10_8,ip_10_9,ip_10_10,ip_10_11,ip_10_12,ip_10_13,ip_10_14,ip_10_15,ip_10_16,ip_10_17,ip_10_18,ip_10_19,ip_10_20,ip_10_21,ip_10_22,ip_10_23,ip_10_24,ip_10_25,ip_10_26,ip_10_27,ip_10_28,ip_10_29,ip_10_30,ip_10_31,ip_10_32,ip_10_33,ip_10_34,ip_10_35,ip_10_36,ip_10_37,ip_10_38,ip_10_39,ip_10_40,ip_10_41,ip_10_42,ip_10_43,ip_10_44,ip_10_45,ip_10_46,ip_10_47,ip_10_48,ip_10_49,ip_10_50,ip_10_51,ip_10_52,ip_10_53,ip_10_54,ip_10_55,ip_10_56,ip_10_57,ip_10_58,ip_10_59,ip_10_60,ip_10_61,ip_10_62,ip_10_63,ip_11_0,ip_11_1,ip_11_2,ip_11_3,ip_11_4,ip_11_5,ip_11_6,ip_11_7,ip_11_8,ip_11_9,ip_11_10,ip_11_11,ip_11_12,ip_11_13,ip_11_14,ip_11_15,ip_11_16,ip_11_17,ip_11_18,ip_11_19,ip_11_20,ip_11_21,ip_11_22,ip_11_23,ip_11_24,ip_11_25,ip_11_26,ip_11_27,ip_11_28,ip_11_29,ip_11_30,ip_11_31,ip_11_32,ip_11_33,ip_11_34,ip_11_35,ip_11_36,ip_11_37,ip_11_38,ip_11_39,ip_11_40,ip_11_41,ip_11_42,ip_11_43,ip_11_44,ip_11_45,ip_11_46,ip_11_47,ip_11_48,ip_11_49,ip_11_50,ip_11_51,ip_11_52,ip_11_53,ip_11_54,ip_11_55,ip_11_56,ip_11_57,ip_11_58,ip_11_59,ip_11_60,ip_11_61,ip_11_62,ip_11_63,ip_12_0,ip_12_1,ip_12_2,ip_12_3,ip_12_4,ip_12_5,ip_12_6,ip_12_7,ip_12_8,ip_12_9,ip_12_10,ip_12_11,ip_12_12,ip_12_13,ip_12_14,ip_12_15,ip_12_16,ip_12_17,ip_12_18,ip_12_19,ip_12_20,ip_12_21,ip_12_22,ip_12_23,ip_12_24,ip_12_25,ip_12_26,ip_12_27,ip_12_28,ip_12_29,ip_12_30,ip_12_31,ip_12_32,ip_12_33,ip_12_34,ip_12_35,ip_12_36,ip_12_37,ip_12_38,ip_12_39,ip_12_40,ip_12_41,ip_12_42,ip_12_43,ip_12_44,ip_12_45,ip_12_46,ip_12_47,ip_12_48,ip_12_49,ip_12_50,ip_12_51,ip_12_52,ip_12_53,ip_12_54,ip_12_55,ip_12_56,ip_12_57,ip_12_58,ip_12_59,ip_12_60,ip_12_61,ip_12_62,ip_12_63,ip_13_0,ip_13_1,ip_13_2,ip_13_3,ip_13_4,ip_13_5,ip_13_6,ip_13_7,ip_13_8,ip_13_9,ip_13_10,ip_13_11,ip_13_12,ip_13_13,ip_13_14,ip_13_15,ip_13_16,ip_13_17,ip_13_18,ip_13_19,ip_13_20,ip_13_21,ip_13_22,ip_13_23,ip_13_24,ip_13_25,ip_13_26,ip_13_27,ip_13_28,ip_13_29,ip_13_30,ip_13_31,ip_13_32,ip_13_33,ip_13_34,ip_13_35,ip_13_36,ip_13_37,ip_13_38,ip_13_39,ip_13_40,ip_13_41,ip_13_42,ip_13_43,ip_13_44,ip_13_45,ip_13_46,ip_13_47,ip_13_48,ip_13_49,ip_13_50,ip_13_51,ip_13_52,ip_13_53,ip_13_54,ip_13_55,ip_13_56,ip_13_57,ip_13_58,ip_13_59,ip_13_60,ip_13_61,ip_13_62,ip_13_63,ip_14_0,ip_14_1,ip_14_2,ip_14_3,ip_14_4,ip_14_5,ip_14_6,ip_14_7,ip_14_8,ip_14_9,ip_14_10,ip_14_11,ip_14_12,ip_14_13,ip_14_14,ip_14_15,ip_14_16,ip_14_17,ip_14_18,ip_14_19,ip_14_20,ip_14_21,ip_14_22,ip_14_23,ip_14_24,ip_14_25,ip_14_26,ip_14_27,ip_14_28,ip_14_29,ip_14_30,ip_14_31,ip_14_32,ip_14_33,ip_14_34,ip_14_35,ip_14_36,ip_14_37,ip_14_38,ip_14_39,ip_14_40,ip_14_41,ip_14_42,ip_14_43,ip_14_44,ip_14_45,ip_14_46,ip_14_47,ip_14_48,ip_14_49,ip_14_50,ip_14_51,ip_14_52,ip_14_53,ip_14_54,ip_14_55,ip_14_56,ip_14_57,ip_14_58,ip_14_59,ip_14_60,ip_14_61,ip_14_62,ip_14_63,ip_15_0,ip_15_1,ip_15_2,ip_15_3,ip_15_4,ip_15_5,ip_15_6,ip_15_7,ip_15_8,ip_15_9,ip_15_10,ip_15_11,ip_15_12,ip_15_13,ip_15_14,ip_15_15,ip_15_16,ip_15_17,ip_15_18,ip_15_19,ip_15_20,ip_15_21,ip_15_22,ip_15_23,ip_15_24,ip_15_25,ip_15_26,ip_15_27,ip_15_28,ip_15_29,ip_15_30,ip_15_31,ip_15_32,ip_15_33,ip_15_34,ip_15_35,ip_15_36,ip_15_37,ip_15_38,ip_15_39,ip_15_40,ip_15_41,ip_15_42,ip_15_43,ip_15_44,ip_15_45,ip_15_46,ip_15_47,ip_15_48,ip_15_49,ip_15_50,ip_15_51,ip_15_52,ip_15_53,ip_15_54,ip_15_55,ip_15_56,ip_15_57,ip_15_58,ip_15_59,ip_15_60,ip_15_61,ip_15_62,ip_15_63,ip_16_0,ip_16_1,ip_16_2,ip_16_3,ip_16_4,ip_16_5,ip_16_6,ip_16_7,ip_16_8,ip_16_9,ip_16_10,ip_16_11,ip_16_12,ip_16_13,ip_16_14,ip_16_15,ip_16_16,ip_16_17,ip_16_18,ip_16_19,ip_16_20,ip_16_21,ip_16_22,ip_16_23,ip_16_24,ip_16_25,ip_16_26,ip_16_27,ip_16_28,ip_16_29,ip_16_30,ip_16_31,ip_16_32,ip_16_33,ip_16_34,ip_16_35,ip_16_36,ip_16_37,ip_16_38,ip_16_39,ip_16_40,ip_16_41,ip_16_42,ip_16_43,ip_16_44,ip_16_45,ip_16_46,ip_16_47,ip_16_48,ip_16_49,ip_16_50,ip_16_51,ip_16_52,ip_16_53,ip_16_54,ip_16_55,ip_16_56,ip_16_57,ip_16_58,ip_16_59,ip_16_60,ip_16_61,ip_16_62,ip_16_63,ip_17_0,ip_17_1,ip_17_2,ip_17_3,ip_17_4,ip_17_5,ip_17_6,ip_17_7,ip_17_8,ip_17_9,ip_17_10,ip_17_11,ip_17_12,ip_17_13,ip_17_14,ip_17_15,ip_17_16,ip_17_17,ip_17_18,ip_17_19,ip_17_20,ip_17_21,ip_17_22,ip_17_23,ip_17_24,ip_17_25,ip_17_26,ip_17_27,ip_17_28,ip_17_29,ip_17_30,ip_17_31,ip_17_32,ip_17_33,ip_17_34,ip_17_35,ip_17_36,ip_17_37,ip_17_38,ip_17_39,ip_17_40,ip_17_41,ip_17_42,ip_17_43,ip_17_44,ip_17_45,ip_17_46,ip_17_47,ip_17_48,ip_17_49,ip_17_50,ip_17_51,ip_17_52,ip_17_53,ip_17_54,ip_17_55,ip_17_56,ip_17_57,ip_17_58,ip_17_59,ip_17_60,ip_17_61,ip_17_62,ip_17_63,ip_18_0,ip_18_1,ip_18_2,ip_18_3,ip_18_4,ip_18_5,ip_18_6,ip_18_7,ip_18_8,ip_18_9,ip_18_10,ip_18_11,ip_18_12,ip_18_13,ip_18_14,ip_18_15,ip_18_16,ip_18_17,ip_18_18,ip_18_19,ip_18_20,ip_18_21,ip_18_22,ip_18_23,ip_18_24,ip_18_25,ip_18_26,ip_18_27,ip_18_28,ip_18_29,ip_18_30,ip_18_31,ip_18_32,ip_18_33,ip_18_34,ip_18_35,ip_18_36,ip_18_37,ip_18_38,ip_18_39,ip_18_40,ip_18_41,ip_18_42,ip_18_43,ip_18_44,ip_18_45,ip_18_46,ip_18_47,ip_18_48,ip_18_49,ip_18_50,ip_18_51,ip_18_52,ip_18_53,ip_18_54,ip_18_55,ip_18_56,ip_18_57,ip_18_58,ip_18_59,ip_18_60,ip_18_61,ip_18_62,ip_18_63,ip_19_0,ip_19_1,ip_19_2,ip_19_3,ip_19_4,ip_19_5,ip_19_6,ip_19_7,ip_19_8,ip_19_9,ip_19_10,ip_19_11,ip_19_12,ip_19_13,ip_19_14,ip_19_15,ip_19_16,ip_19_17,ip_19_18,ip_19_19,ip_19_20,ip_19_21,ip_19_22,ip_19_23,ip_19_24,ip_19_25,ip_19_26,ip_19_27,ip_19_28,ip_19_29,ip_19_30,ip_19_31,ip_19_32,ip_19_33,ip_19_34,ip_19_35,ip_19_36,ip_19_37,ip_19_38,ip_19_39,ip_19_40,ip_19_41,ip_19_42,ip_19_43,ip_19_44,ip_19_45,ip_19_46,ip_19_47,ip_19_48,ip_19_49,ip_19_50,ip_19_51,ip_19_52,ip_19_53,ip_19_54,ip_19_55,ip_19_56,ip_19_57,ip_19_58,ip_19_59,ip_19_60,ip_19_61,ip_19_62,ip_19_63,ip_20_0,ip_20_1,ip_20_2,ip_20_3,ip_20_4,ip_20_5,ip_20_6,ip_20_7,ip_20_8,ip_20_9,ip_20_10,ip_20_11,ip_20_12,ip_20_13,ip_20_14,ip_20_15,ip_20_16,ip_20_17,ip_20_18,ip_20_19,ip_20_20,ip_20_21,ip_20_22,ip_20_23,ip_20_24,ip_20_25,ip_20_26,ip_20_27,ip_20_28,ip_20_29,ip_20_30,ip_20_31,ip_20_32,ip_20_33,ip_20_34,ip_20_35,ip_20_36,ip_20_37,ip_20_38,ip_20_39,ip_20_40,ip_20_41,ip_20_42,ip_20_43,ip_20_44,ip_20_45,ip_20_46,ip_20_47,ip_20_48,ip_20_49,ip_20_50,ip_20_51,ip_20_52,ip_20_53,ip_20_54,ip_20_55,ip_20_56,ip_20_57,ip_20_58,ip_20_59,ip_20_60,ip_20_61,ip_20_62,ip_20_63,ip_21_0,ip_21_1,ip_21_2,ip_21_3,ip_21_4,ip_21_5,ip_21_6,ip_21_7,ip_21_8,ip_21_9,ip_21_10,ip_21_11,ip_21_12,ip_21_13,ip_21_14,ip_21_15,ip_21_16,ip_21_17,ip_21_18,ip_21_19,ip_21_20,ip_21_21,ip_21_22,ip_21_23,ip_21_24,ip_21_25,ip_21_26,ip_21_27,ip_21_28,ip_21_29,ip_21_30,ip_21_31,ip_21_32,ip_21_33,ip_21_34,ip_21_35,ip_21_36,ip_21_37,ip_21_38,ip_21_39,ip_21_40,ip_21_41,ip_21_42,ip_21_43,ip_21_44,ip_21_45,ip_21_46,ip_21_47,ip_21_48,ip_21_49,ip_21_50,ip_21_51,ip_21_52,ip_21_53,ip_21_54,ip_21_55,ip_21_56,ip_21_57,ip_21_58,ip_21_59,ip_21_60,ip_21_61,ip_21_62,ip_21_63,ip_22_0,ip_22_1,ip_22_2,ip_22_3,ip_22_4,ip_22_5,ip_22_6,ip_22_7,ip_22_8,ip_22_9,ip_22_10,ip_22_11,ip_22_12,ip_22_13,ip_22_14,ip_22_15,ip_22_16,ip_22_17,ip_22_18,ip_22_19,ip_22_20,ip_22_21,ip_22_22,ip_22_23,ip_22_24,ip_22_25,ip_22_26,ip_22_27,ip_22_28,ip_22_29,ip_22_30,ip_22_31,ip_22_32,ip_22_33,ip_22_34,ip_22_35,ip_22_36,ip_22_37,ip_22_38,ip_22_39,ip_22_40,ip_22_41,ip_22_42,ip_22_43,ip_22_44,ip_22_45,ip_22_46,ip_22_47,ip_22_48,ip_22_49,ip_22_50,ip_22_51,ip_22_52,ip_22_53,ip_22_54,ip_22_55,ip_22_56,ip_22_57,ip_22_58,ip_22_59,ip_22_60,ip_22_61,ip_22_62,ip_22_63,ip_23_0,ip_23_1,ip_23_2,ip_23_3,ip_23_4,ip_23_5,ip_23_6,ip_23_7,ip_23_8,ip_23_9,ip_23_10,ip_23_11,ip_23_12,ip_23_13,ip_23_14,ip_23_15,ip_23_16,ip_23_17,ip_23_18,ip_23_19,ip_23_20,ip_23_21,ip_23_22,ip_23_23,ip_23_24,ip_23_25,ip_23_26,ip_23_27,ip_23_28,ip_23_29,ip_23_30,ip_23_31,ip_23_32,ip_23_33,ip_23_34,ip_23_35,ip_23_36,ip_23_37,ip_23_38,ip_23_39,ip_23_40,ip_23_41,ip_23_42,ip_23_43,ip_23_44,ip_23_45,ip_23_46,ip_23_47,ip_23_48,ip_23_49,ip_23_50,ip_23_51,ip_23_52,ip_23_53,ip_23_54,ip_23_55,ip_23_56,ip_23_57,ip_23_58,ip_23_59,ip_23_60,ip_23_61,ip_23_62,ip_23_63,ip_24_0,ip_24_1,ip_24_2,ip_24_3,ip_24_4,ip_24_5,ip_24_6,ip_24_7,ip_24_8,ip_24_9,ip_24_10,ip_24_11,ip_24_12,ip_24_13,ip_24_14,ip_24_15,ip_24_16,ip_24_17,ip_24_18,ip_24_19,ip_24_20,ip_24_21,ip_24_22,ip_24_23,ip_24_24,ip_24_25,ip_24_26,ip_24_27,ip_24_28,ip_24_29,ip_24_30,ip_24_31,ip_24_32,ip_24_33,ip_24_34,ip_24_35,ip_24_36,ip_24_37,ip_24_38,ip_24_39,ip_24_40,ip_24_41,ip_24_42,ip_24_43,ip_24_44,ip_24_45,ip_24_46,ip_24_47,ip_24_48,ip_24_49,ip_24_50,ip_24_51,ip_24_52,ip_24_53,ip_24_54,ip_24_55,ip_24_56,ip_24_57,ip_24_58,ip_24_59,ip_24_60,ip_24_61,ip_24_62,ip_24_63,ip_25_0,ip_25_1,ip_25_2,ip_25_3,ip_25_4,ip_25_5,ip_25_6,ip_25_7,ip_25_8,ip_25_9,ip_25_10,ip_25_11,ip_25_12,ip_25_13,ip_25_14,ip_25_15,ip_25_16,ip_25_17,ip_25_18,ip_25_19,ip_25_20,ip_25_21,ip_25_22,ip_25_23,ip_25_24,ip_25_25,ip_25_26,ip_25_27,ip_25_28,ip_25_29,ip_25_30,ip_25_31,ip_25_32,ip_25_33,ip_25_34,ip_25_35,ip_25_36,ip_25_37,ip_25_38,ip_25_39,ip_25_40,ip_25_41,ip_25_42,ip_25_43,ip_25_44,ip_25_45,ip_25_46,ip_25_47,ip_25_48,ip_25_49,ip_25_50,ip_25_51,ip_25_52,ip_25_53,ip_25_54,ip_25_55,ip_25_56,ip_25_57,ip_25_58,ip_25_59,ip_25_60,ip_25_61,ip_25_62,ip_25_63,ip_26_0,ip_26_1,ip_26_2,ip_26_3,ip_26_4,ip_26_5,ip_26_6,ip_26_7,ip_26_8,ip_26_9,ip_26_10,ip_26_11,ip_26_12,ip_26_13,ip_26_14,ip_26_15,ip_26_16,ip_26_17,ip_26_18,ip_26_19,ip_26_20,ip_26_21,ip_26_22,ip_26_23,ip_26_24,ip_26_25,ip_26_26,ip_26_27,ip_26_28,ip_26_29,ip_26_30,ip_26_31,ip_26_32,ip_26_33,ip_26_34,ip_26_35,ip_26_36,ip_26_37,ip_26_38,ip_26_39,ip_26_40,ip_26_41,ip_26_42,ip_26_43,ip_26_44,ip_26_45,ip_26_46,ip_26_47,ip_26_48,ip_26_49,ip_26_50,ip_26_51,ip_26_52,ip_26_53,ip_26_54,ip_26_55,ip_26_56,ip_26_57,ip_26_58,ip_26_59,ip_26_60,ip_26_61,ip_26_62,ip_26_63,ip_27_0,ip_27_1,ip_27_2,ip_27_3,ip_27_4,ip_27_5,ip_27_6,ip_27_7,ip_27_8,ip_27_9,ip_27_10,ip_27_11,ip_27_12,ip_27_13,ip_27_14,ip_27_15,ip_27_16,ip_27_17,ip_27_18,ip_27_19,ip_27_20,ip_27_21,ip_27_22,ip_27_23,ip_27_24,ip_27_25,ip_27_26,ip_27_27,ip_27_28,ip_27_29,ip_27_30,ip_27_31,ip_27_32,ip_27_33,ip_27_34,ip_27_35,ip_27_36,ip_27_37,ip_27_38,ip_27_39,ip_27_40,ip_27_41,ip_27_42,ip_27_43,ip_27_44,ip_27_45,ip_27_46,ip_27_47,ip_27_48,ip_27_49,ip_27_50,ip_27_51,ip_27_52,ip_27_53,ip_27_54,ip_27_55,ip_27_56,ip_27_57,ip_27_58,ip_27_59,ip_27_60,ip_27_61,ip_27_62,ip_27_63,ip_28_0,ip_28_1,ip_28_2,ip_28_3,ip_28_4,ip_28_5,ip_28_6,ip_28_7,ip_28_8,ip_28_9,ip_28_10,ip_28_11,ip_28_12,ip_28_13,ip_28_14,ip_28_15,ip_28_16,ip_28_17,ip_28_18,ip_28_19,ip_28_20,ip_28_21,ip_28_22,ip_28_23,ip_28_24,ip_28_25,ip_28_26,ip_28_27,ip_28_28,ip_28_29,ip_28_30,ip_28_31,ip_28_32,ip_28_33,ip_28_34,ip_28_35,ip_28_36,ip_28_37,ip_28_38,ip_28_39,ip_28_40,ip_28_41,ip_28_42,ip_28_43,ip_28_44,ip_28_45,ip_28_46,ip_28_47,ip_28_48,ip_28_49,ip_28_50,ip_28_51,ip_28_52,ip_28_53,ip_28_54,ip_28_55,ip_28_56,ip_28_57,ip_28_58,ip_28_59,ip_28_60,ip_28_61,ip_28_62,ip_28_63,ip_29_0,ip_29_1,ip_29_2,ip_29_3,ip_29_4,ip_29_5,ip_29_6,ip_29_7,ip_29_8,ip_29_9,ip_29_10,ip_29_11,ip_29_12,ip_29_13,ip_29_14,ip_29_15,ip_29_16,ip_29_17,ip_29_18,ip_29_19,ip_29_20,ip_29_21,ip_29_22,ip_29_23,ip_29_24,ip_29_25,ip_29_26,ip_29_27,ip_29_28,ip_29_29,ip_29_30,ip_29_31,ip_29_32,ip_29_33,ip_29_34,ip_29_35,ip_29_36,ip_29_37,ip_29_38,ip_29_39,ip_29_40,ip_29_41,ip_29_42,ip_29_43,ip_29_44,ip_29_45,ip_29_46,ip_29_47,ip_29_48,ip_29_49,ip_29_50,ip_29_51,ip_29_52,ip_29_53,ip_29_54,ip_29_55,ip_29_56,ip_29_57,ip_29_58,ip_29_59,ip_29_60,ip_29_61,ip_29_62,ip_29_63,ip_30_0,ip_30_1,ip_30_2,ip_30_3,ip_30_4,ip_30_5,ip_30_6,ip_30_7,ip_30_8,ip_30_9,ip_30_10,ip_30_11,ip_30_12,ip_30_13,ip_30_14,ip_30_15,ip_30_16,ip_30_17,ip_30_18,ip_30_19,ip_30_20,ip_30_21,ip_30_22,ip_30_23,ip_30_24,ip_30_25,ip_30_26,ip_30_27,ip_30_28,ip_30_29,ip_30_30,ip_30_31,ip_30_32,ip_30_33,ip_30_34,ip_30_35,ip_30_36,ip_30_37,ip_30_38,ip_30_39,ip_30_40,ip_30_41,ip_30_42,ip_30_43,ip_30_44,ip_30_45,ip_30_46,ip_30_47,ip_30_48,ip_30_49,ip_30_50,ip_30_51,ip_30_52,ip_30_53,ip_30_54,ip_30_55,ip_30_56,ip_30_57,ip_30_58,ip_30_59,ip_30_60,ip_30_61,ip_30_62,ip_30_63,ip_31_0,ip_31_1,ip_31_2,ip_31_3,ip_31_4,ip_31_5,ip_31_6,ip_31_7,ip_31_8,ip_31_9,ip_31_10,ip_31_11,ip_31_12,ip_31_13,ip_31_14,ip_31_15,ip_31_16,ip_31_17,ip_31_18,ip_31_19,ip_31_20,ip_31_21,ip_31_22,ip_31_23,ip_31_24,ip_31_25,ip_31_26,ip_31_27,ip_31_28,ip_31_29,ip_31_30,ip_31_31,ip_31_32,ip_31_33,ip_31_34,ip_31_35,ip_31_36,ip_31_37,ip_31_38,ip_31_39,ip_31_40,ip_31_41,ip_31_42,ip_31_43,ip_31_44,ip_31_45,ip_31_46,ip_31_47,ip_31_48,ip_31_49,ip_31_50,ip_31_51,ip_31_52,ip_31_53,ip_31_54,ip_31_55,ip_31_56,ip_31_57,ip_31_58,ip_31_59,ip_31_60,ip_31_61,ip_31_62,ip_31_63,ip_32_0,ip_32_1,ip_32_2,ip_32_3,ip_32_4,ip_32_5,ip_32_6,ip_32_7,ip_32_8,ip_32_9,ip_32_10,ip_32_11,ip_32_12,ip_32_13,ip_32_14,ip_32_15,ip_32_16,ip_32_17,ip_32_18,ip_32_19,ip_32_20,ip_32_21,ip_32_22,ip_32_23,ip_32_24,ip_32_25,ip_32_26,ip_32_27,ip_32_28,ip_32_29,ip_32_30,ip_32_31,ip_32_32,ip_32_33,ip_32_34,ip_32_35,ip_32_36,ip_32_37,ip_32_38,ip_32_39,ip_32_40,ip_32_41,ip_32_42,ip_32_43,ip_32_44,ip_32_45,ip_32_46,ip_32_47,ip_32_48,ip_32_49,ip_32_50,ip_32_51,ip_32_52,ip_32_53,ip_32_54,ip_32_55,ip_32_56,ip_32_57,ip_32_58,ip_32_59,ip_32_60,ip_32_61,ip_32_62,ip_32_63,ip_33_0,ip_33_1,ip_33_2,ip_33_3,ip_33_4,ip_33_5,ip_33_6,ip_33_7,ip_33_8,ip_33_9,ip_33_10,ip_33_11,ip_33_12,ip_33_13,ip_33_14,ip_33_15,ip_33_16,ip_33_17,ip_33_18,ip_33_19,ip_33_20,ip_33_21,ip_33_22,ip_33_23,ip_33_24,ip_33_25,ip_33_26,ip_33_27,ip_33_28,ip_33_29,ip_33_30,ip_33_31,ip_33_32,ip_33_33,ip_33_34,ip_33_35,ip_33_36,ip_33_37,ip_33_38,ip_33_39,ip_33_40,ip_33_41,ip_33_42,ip_33_43,ip_33_44,ip_33_45,ip_33_46,ip_33_47,ip_33_48,ip_33_49,ip_33_50,ip_33_51,ip_33_52,ip_33_53,ip_33_54,ip_33_55,ip_33_56,ip_33_57,ip_33_58,ip_33_59,ip_33_60,ip_33_61,ip_33_62,ip_33_63,ip_34_0,ip_34_1,ip_34_2,ip_34_3,ip_34_4,ip_34_5,ip_34_6,ip_34_7,ip_34_8,ip_34_9,ip_34_10,ip_34_11,ip_34_12,ip_34_13,ip_34_14,ip_34_15,ip_34_16,ip_34_17,ip_34_18,ip_34_19,ip_34_20,ip_34_21,ip_34_22,ip_34_23,ip_34_24,ip_34_25,ip_34_26,ip_34_27,ip_34_28,ip_34_29,ip_34_30,ip_34_31,ip_34_32,ip_34_33,ip_34_34,ip_34_35,ip_34_36,ip_34_37,ip_34_38,ip_34_39,ip_34_40,ip_34_41,ip_34_42,ip_34_43,ip_34_44,ip_34_45,ip_34_46,ip_34_47,ip_34_48,ip_34_49,ip_34_50,ip_34_51,ip_34_52,ip_34_53,ip_34_54,ip_34_55,ip_34_56,ip_34_57,ip_34_58,ip_34_59,ip_34_60,ip_34_61,ip_34_62,ip_34_63,ip_35_0,ip_35_1,ip_35_2,ip_35_3,ip_35_4,ip_35_5,ip_35_6,ip_35_7,ip_35_8,ip_35_9,ip_35_10,ip_35_11,ip_35_12,ip_35_13,ip_35_14,ip_35_15,ip_35_16,ip_35_17,ip_35_18,ip_35_19,ip_35_20,ip_35_21,ip_35_22,ip_35_23,ip_35_24,ip_35_25,ip_35_26,ip_35_27,ip_35_28,ip_35_29,ip_35_30,ip_35_31,ip_35_32,ip_35_33,ip_35_34,ip_35_35,ip_35_36,ip_35_37,ip_35_38,ip_35_39,ip_35_40,ip_35_41,ip_35_42,ip_35_43,ip_35_44,ip_35_45,ip_35_46,ip_35_47,ip_35_48,ip_35_49,ip_35_50,ip_35_51,ip_35_52,ip_35_53,ip_35_54,ip_35_55,ip_35_56,ip_35_57,ip_35_58,ip_35_59,ip_35_60,ip_35_61,ip_35_62,ip_35_63,ip_36_0,ip_36_1,ip_36_2,ip_36_3,ip_36_4,ip_36_5,ip_36_6,ip_36_7,ip_36_8,ip_36_9,ip_36_10,ip_36_11,ip_36_12,ip_36_13,ip_36_14,ip_36_15,ip_36_16,ip_36_17,ip_36_18,ip_36_19,ip_36_20,ip_36_21,ip_36_22,ip_36_23,ip_36_24,ip_36_25,ip_36_26,ip_36_27,ip_36_28,ip_36_29,ip_36_30,ip_36_31,ip_36_32,ip_36_33,ip_36_34,ip_36_35,ip_36_36,ip_36_37,ip_36_38,ip_36_39,ip_36_40,ip_36_41,ip_36_42,ip_36_43,ip_36_44,ip_36_45,ip_36_46,ip_36_47,ip_36_48,ip_36_49,ip_36_50,ip_36_51,ip_36_52,ip_36_53,ip_36_54,ip_36_55,ip_36_56,ip_36_57,ip_36_58,ip_36_59,ip_36_60,ip_36_61,ip_36_62,ip_36_63,ip_37_0,ip_37_1,ip_37_2,ip_37_3,ip_37_4,ip_37_5,ip_37_6,ip_37_7,ip_37_8,ip_37_9,ip_37_10,ip_37_11,ip_37_12,ip_37_13,ip_37_14,ip_37_15,ip_37_16,ip_37_17,ip_37_18,ip_37_19,ip_37_20,ip_37_21,ip_37_22,ip_37_23,ip_37_24,ip_37_25,ip_37_26,ip_37_27,ip_37_28,ip_37_29,ip_37_30,ip_37_31,ip_37_32,ip_37_33,ip_37_34,ip_37_35,ip_37_36,ip_37_37,ip_37_38,ip_37_39,ip_37_40,ip_37_41,ip_37_42,ip_37_43,ip_37_44,ip_37_45,ip_37_46,ip_37_47,ip_37_48,ip_37_49,ip_37_50,ip_37_51,ip_37_52,ip_37_53,ip_37_54,ip_37_55,ip_37_56,ip_37_57,ip_37_58,ip_37_59,ip_37_60,ip_37_61,ip_37_62,ip_37_63,ip_38_0,ip_38_1,ip_38_2,ip_38_3,ip_38_4,ip_38_5,ip_38_6,ip_38_7,ip_38_8,ip_38_9,ip_38_10,ip_38_11,ip_38_12,ip_38_13,ip_38_14,ip_38_15,ip_38_16,ip_38_17,ip_38_18,ip_38_19,ip_38_20,ip_38_21,ip_38_22,ip_38_23,ip_38_24,ip_38_25,ip_38_26,ip_38_27,ip_38_28,ip_38_29,ip_38_30,ip_38_31,ip_38_32,ip_38_33,ip_38_34,ip_38_35,ip_38_36,ip_38_37,ip_38_38,ip_38_39,ip_38_40,ip_38_41,ip_38_42,ip_38_43,ip_38_44,ip_38_45,ip_38_46,ip_38_47,ip_38_48,ip_38_49,ip_38_50,ip_38_51,ip_38_52,ip_38_53,ip_38_54,ip_38_55,ip_38_56,ip_38_57,ip_38_58,ip_38_59,ip_38_60,ip_38_61,ip_38_62,ip_38_63,ip_39_0,ip_39_1,ip_39_2,ip_39_3,ip_39_4,ip_39_5,ip_39_6,ip_39_7,ip_39_8,ip_39_9,ip_39_10,ip_39_11,ip_39_12,ip_39_13,ip_39_14,ip_39_15,ip_39_16,ip_39_17,ip_39_18,ip_39_19,ip_39_20,ip_39_21,ip_39_22,ip_39_23,ip_39_24,ip_39_25,ip_39_26,ip_39_27,ip_39_28,ip_39_29,ip_39_30,ip_39_31,ip_39_32,ip_39_33,ip_39_34,ip_39_35,ip_39_36,ip_39_37,ip_39_38,ip_39_39,ip_39_40,ip_39_41,ip_39_42,ip_39_43,ip_39_44,ip_39_45,ip_39_46,ip_39_47,ip_39_48,ip_39_49,ip_39_50,ip_39_51,ip_39_52,ip_39_53,ip_39_54,ip_39_55,ip_39_56,ip_39_57,ip_39_58,ip_39_59,ip_39_60,ip_39_61,ip_39_62,ip_39_63,ip_40_0,ip_40_1,ip_40_2,ip_40_3,ip_40_4,ip_40_5,ip_40_6,ip_40_7,ip_40_8,ip_40_9,ip_40_10,ip_40_11,ip_40_12,ip_40_13,ip_40_14,ip_40_15,ip_40_16,ip_40_17,ip_40_18,ip_40_19,ip_40_20,ip_40_21,ip_40_22,ip_40_23,ip_40_24,ip_40_25,ip_40_26,ip_40_27,ip_40_28,ip_40_29,ip_40_30,ip_40_31,ip_40_32,ip_40_33,ip_40_34,ip_40_35,ip_40_36,ip_40_37,ip_40_38,ip_40_39,ip_40_40,ip_40_41,ip_40_42,ip_40_43,ip_40_44,ip_40_45,ip_40_46,ip_40_47,ip_40_48,ip_40_49,ip_40_50,ip_40_51,ip_40_52,ip_40_53,ip_40_54,ip_40_55,ip_40_56,ip_40_57,ip_40_58,ip_40_59,ip_40_60,ip_40_61,ip_40_62,ip_40_63,ip_41_0,ip_41_1,ip_41_2,ip_41_3,ip_41_4,ip_41_5,ip_41_6,ip_41_7,ip_41_8,ip_41_9,ip_41_10,ip_41_11,ip_41_12,ip_41_13,ip_41_14,ip_41_15,ip_41_16,ip_41_17,ip_41_18,ip_41_19,ip_41_20,ip_41_21,ip_41_22,ip_41_23,ip_41_24,ip_41_25,ip_41_26,ip_41_27,ip_41_28,ip_41_29,ip_41_30,ip_41_31,ip_41_32,ip_41_33,ip_41_34,ip_41_35,ip_41_36,ip_41_37,ip_41_38,ip_41_39,ip_41_40,ip_41_41,ip_41_42,ip_41_43,ip_41_44,ip_41_45,ip_41_46,ip_41_47,ip_41_48,ip_41_49,ip_41_50,ip_41_51,ip_41_52,ip_41_53,ip_41_54,ip_41_55,ip_41_56,ip_41_57,ip_41_58,ip_41_59,ip_41_60,ip_41_61,ip_41_62,ip_41_63,ip_42_0,ip_42_1,ip_42_2,ip_42_3,ip_42_4,ip_42_5,ip_42_6,ip_42_7,ip_42_8,ip_42_9,ip_42_10,ip_42_11,ip_42_12,ip_42_13,ip_42_14,ip_42_15,ip_42_16,ip_42_17,ip_42_18,ip_42_19,ip_42_20,ip_42_21,ip_42_22,ip_42_23,ip_42_24,ip_42_25,ip_42_26,ip_42_27,ip_42_28,ip_42_29,ip_42_30,ip_42_31,ip_42_32,ip_42_33,ip_42_34,ip_42_35,ip_42_36,ip_42_37,ip_42_38,ip_42_39,ip_42_40,ip_42_41,ip_42_42,ip_42_43,ip_42_44,ip_42_45,ip_42_46,ip_42_47,ip_42_48,ip_42_49,ip_42_50,ip_42_51,ip_42_52,ip_42_53,ip_42_54,ip_42_55,ip_42_56,ip_42_57,ip_42_58,ip_42_59,ip_42_60,ip_42_61,ip_42_62,ip_42_63,ip_43_0,ip_43_1,ip_43_2,ip_43_3,ip_43_4,ip_43_5,ip_43_6,ip_43_7,ip_43_8,ip_43_9,ip_43_10,ip_43_11,ip_43_12,ip_43_13,ip_43_14,ip_43_15,ip_43_16,ip_43_17,ip_43_18,ip_43_19,ip_43_20,ip_43_21,ip_43_22,ip_43_23,ip_43_24,ip_43_25,ip_43_26,ip_43_27,ip_43_28,ip_43_29,ip_43_30,ip_43_31,ip_43_32,ip_43_33,ip_43_34,ip_43_35,ip_43_36,ip_43_37,ip_43_38,ip_43_39,ip_43_40,ip_43_41,ip_43_42,ip_43_43,ip_43_44,ip_43_45,ip_43_46,ip_43_47,ip_43_48,ip_43_49,ip_43_50,ip_43_51,ip_43_52,ip_43_53,ip_43_54,ip_43_55,ip_43_56,ip_43_57,ip_43_58,ip_43_59,ip_43_60,ip_43_61,ip_43_62,ip_43_63,ip_44_0,ip_44_1,ip_44_2,ip_44_3,ip_44_4,ip_44_5,ip_44_6,ip_44_7,ip_44_8,ip_44_9,ip_44_10,ip_44_11,ip_44_12,ip_44_13,ip_44_14,ip_44_15,ip_44_16,ip_44_17,ip_44_18,ip_44_19,ip_44_20,ip_44_21,ip_44_22,ip_44_23,ip_44_24,ip_44_25,ip_44_26,ip_44_27,ip_44_28,ip_44_29,ip_44_30,ip_44_31,ip_44_32,ip_44_33,ip_44_34,ip_44_35,ip_44_36,ip_44_37,ip_44_38,ip_44_39,ip_44_40,ip_44_41,ip_44_42,ip_44_43,ip_44_44,ip_44_45,ip_44_46,ip_44_47,ip_44_48,ip_44_49,ip_44_50,ip_44_51,ip_44_52,ip_44_53,ip_44_54,ip_44_55,ip_44_56,ip_44_57,ip_44_58,ip_44_59,ip_44_60,ip_44_61,ip_44_62,ip_44_63,ip_45_0,ip_45_1,ip_45_2,ip_45_3,ip_45_4,ip_45_5,ip_45_6,ip_45_7,ip_45_8,ip_45_9,ip_45_10,ip_45_11,ip_45_12,ip_45_13,ip_45_14,ip_45_15,ip_45_16,ip_45_17,ip_45_18,ip_45_19,ip_45_20,ip_45_21,ip_45_22,ip_45_23,ip_45_24,ip_45_25,ip_45_26,ip_45_27,ip_45_28,ip_45_29,ip_45_30,ip_45_31,ip_45_32,ip_45_33,ip_45_34,ip_45_35,ip_45_36,ip_45_37,ip_45_38,ip_45_39,ip_45_40,ip_45_41,ip_45_42,ip_45_43,ip_45_44,ip_45_45,ip_45_46,ip_45_47,ip_45_48,ip_45_49,ip_45_50,ip_45_51,ip_45_52,ip_45_53,ip_45_54,ip_45_55,ip_45_56,ip_45_57,ip_45_58,ip_45_59,ip_45_60,ip_45_61,ip_45_62,ip_45_63,ip_46_0,ip_46_1,ip_46_2,ip_46_3,ip_46_4,ip_46_5,ip_46_6,ip_46_7,ip_46_8,ip_46_9,ip_46_10,ip_46_11,ip_46_12,ip_46_13,ip_46_14,ip_46_15,ip_46_16,ip_46_17,ip_46_18,ip_46_19,ip_46_20,ip_46_21,ip_46_22,ip_46_23,ip_46_24,ip_46_25,ip_46_26,ip_46_27,ip_46_28,ip_46_29,ip_46_30,ip_46_31,ip_46_32,ip_46_33,ip_46_34,ip_46_35,ip_46_36,ip_46_37,ip_46_38,ip_46_39,ip_46_40,ip_46_41,ip_46_42,ip_46_43,ip_46_44,ip_46_45,ip_46_46,ip_46_47,ip_46_48,ip_46_49,ip_46_50,ip_46_51,ip_46_52,ip_46_53,ip_46_54,ip_46_55,ip_46_56,ip_46_57,ip_46_58,ip_46_59,ip_46_60,ip_46_61,ip_46_62,ip_46_63,ip_47_0,ip_47_1,ip_47_2,ip_47_3,ip_47_4,ip_47_5,ip_47_6,ip_47_7,ip_47_8,ip_47_9,ip_47_10,ip_47_11,ip_47_12,ip_47_13,ip_47_14,ip_47_15,ip_47_16,ip_47_17,ip_47_18,ip_47_19,ip_47_20,ip_47_21,ip_47_22,ip_47_23,ip_47_24,ip_47_25,ip_47_26,ip_47_27,ip_47_28,ip_47_29,ip_47_30,ip_47_31,ip_47_32,ip_47_33,ip_47_34,ip_47_35,ip_47_36,ip_47_37,ip_47_38,ip_47_39,ip_47_40,ip_47_41,ip_47_42,ip_47_43,ip_47_44,ip_47_45,ip_47_46,ip_47_47,ip_47_48,ip_47_49,ip_47_50,ip_47_51,ip_47_52,ip_47_53,ip_47_54,ip_47_55,ip_47_56,ip_47_57,ip_47_58,ip_47_59,ip_47_60,ip_47_61,ip_47_62,ip_47_63,ip_48_0,ip_48_1,ip_48_2,ip_48_3,ip_48_4,ip_48_5,ip_48_6,ip_48_7,ip_48_8,ip_48_9,ip_48_10,ip_48_11,ip_48_12,ip_48_13,ip_48_14,ip_48_15,ip_48_16,ip_48_17,ip_48_18,ip_48_19,ip_48_20,ip_48_21,ip_48_22,ip_48_23,ip_48_24,ip_48_25,ip_48_26,ip_48_27,ip_48_28,ip_48_29,ip_48_30,ip_48_31,ip_48_32,ip_48_33,ip_48_34,ip_48_35,ip_48_36,ip_48_37,ip_48_38,ip_48_39,ip_48_40,ip_48_41,ip_48_42,ip_48_43,ip_48_44,ip_48_45,ip_48_46,ip_48_47,ip_48_48,ip_48_49,ip_48_50,ip_48_51,ip_48_52,ip_48_53,ip_48_54,ip_48_55,ip_48_56,ip_48_57,ip_48_58,ip_48_59,ip_48_60,ip_48_61,ip_48_62,ip_48_63,ip_49_0,ip_49_1,ip_49_2,ip_49_3,ip_49_4,ip_49_5,ip_49_6,ip_49_7,ip_49_8,ip_49_9,ip_49_10,ip_49_11,ip_49_12,ip_49_13,ip_49_14,ip_49_15,ip_49_16,ip_49_17,ip_49_18,ip_49_19,ip_49_20,ip_49_21,ip_49_22,ip_49_23,ip_49_24,ip_49_25,ip_49_26,ip_49_27,ip_49_28,ip_49_29,ip_49_30,ip_49_31,ip_49_32,ip_49_33,ip_49_34,ip_49_35,ip_49_36,ip_49_37,ip_49_38,ip_49_39,ip_49_40,ip_49_41,ip_49_42,ip_49_43,ip_49_44,ip_49_45,ip_49_46,ip_49_47,ip_49_48,ip_49_49,ip_49_50,ip_49_51,ip_49_52,ip_49_53,ip_49_54,ip_49_55,ip_49_56,ip_49_57,ip_49_58,ip_49_59,ip_49_60,ip_49_61,ip_49_62,ip_49_63,ip_50_0,ip_50_1,ip_50_2,ip_50_3,ip_50_4,ip_50_5,ip_50_6,ip_50_7,ip_50_8,ip_50_9,ip_50_10,ip_50_11,ip_50_12,ip_50_13,ip_50_14,ip_50_15,ip_50_16,ip_50_17,ip_50_18,ip_50_19,ip_50_20,ip_50_21,ip_50_22,ip_50_23,ip_50_24,ip_50_25,ip_50_26,ip_50_27,ip_50_28,ip_50_29,ip_50_30,ip_50_31,ip_50_32,ip_50_33,ip_50_34,ip_50_35,ip_50_36,ip_50_37,ip_50_38,ip_50_39,ip_50_40,ip_50_41,ip_50_42,ip_50_43,ip_50_44,ip_50_45,ip_50_46,ip_50_47,ip_50_48,ip_50_49,ip_50_50,ip_50_51,ip_50_52,ip_50_53,ip_50_54,ip_50_55,ip_50_56,ip_50_57,ip_50_58,ip_50_59,ip_50_60,ip_50_61,ip_50_62,ip_50_63,ip_51_0,ip_51_1,ip_51_2,ip_51_3,ip_51_4,ip_51_5,ip_51_6,ip_51_7,ip_51_8,ip_51_9,ip_51_10,ip_51_11,ip_51_12,ip_51_13,ip_51_14,ip_51_15,ip_51_16,ip_51_17,ip_51_18,ip_51_19,ip_51_20,ip_51_21,ip_51_22,ip_51_23,ip_51_24,ip_51_25,ip_51_26,ip_51_27,ip_51_28,ip_51_29,ip_51_30,ip_51_31,ip_51_32,ip_51_33,ip_51_34,ip_51_35,ip_51_36,ip_51_37,ip_51_38,ip_51_39,ip_51_40,ip_51_41,ip_51_42,ip_51_43,ip_51_44,ip_51_45,ip_51_46,ip_51_47,ip_51_48,ip_51_49,ip_51_50,ip_51_51,ip_51_52,ip_51_53,ip_51_54,ip_51_55,ip_51_56,ip_51_57,ip_51_58,ip_51_59,ip_51_60,ip_51_61,ip_51_62,ip_51_63,ip_52_0,ip_52_1,ip_52_2,ip_52_3,ip_52_4,ip_52_5,ip_52_6,ip_52_7,ip_52_8,ip_52_9,ip_52_10,ip_52_11,ip_52_12,ip_52_13,ip_52_14,ip_52_15,ip_52_16,ip_52_17,ip_52_18,ip_52_19,ip_52_20,ip_52_21,ip_52_22,ip_52_23,ip_52_24,ip_52_25,ip_52_26,ip_52_27,ip_52_28,ip_52_29,ip_52_30,ip_52_31,ip_52_32,ip_52_33,ip_52_34,ip_52_35,ip_52_36,ip_52_37,ip_52_38,ip_52_39,ip_52_40,ip_52_41,ip_52_42,ip_52_43,ip_52_44,ip_52_45,ip_52_46,ip_52_47,ip_52_48,ip_52_49,ip_52_50,ip_52_51,ip_52_52,ip_52_53,ip_52_54,ip_52_55,ip_52_56,ip_52_57,ip_52_58,ip_52_59,ip_52_60,ip_52_61,ip_52_62,ip_52_63,ip_53_0,ip_53_1,ip_53_2,ip_53_3,ip_53_4,ip_53_5,ip_53_6,ip_53_7,ip_53_8,ip_53_9,ip_53_10,ip_53_11,ip_53_12,ip_53_13,ip_53_14,ip_53_15,ip_53_16,ip_53_17,ip_53_18,ip_53_19,ip_53_20,ip_53_21,ip_53_22,ip_53_23,ip_53_24,ip_53_25,ip_53_26,ip_53_27,ip_53_28,ip_53_29,ip_53_30,ip_53_31,ip_53_32,ip_53_33,ip_53_34,ip_53_35,ip_53_36,ip_53_37,ip_53_38,ip_53_39,ip_53_40,ip_53_41,ip_53_42,ip_53_43,ip_53_44,ip_53_45,ip_53_46,ip_53_47,ip_53_48,ip_53_49,ip_53_50,ip_53_51,ip_53_52,ip_53_53,ip_53_54,ip_53_55,ip_53_56,ip_53_57,ip_53_58,ip_53_59,ip_53_60,ip_53_61,ip_53_62,ip_53_63,ip_54_0,ip_54_1,ip_54_2,ip_54_3,ip_54_4,ip_54_5,ip_54_6,ip_54_7,ip_54_8,ip_54_9,ip_54_10,ip_54_11,ip_54_12,ip_54_13,ip_54_14,ip_54_15,ip_54_16,ip_54_17,ip_54_18,ip_54_19,ip_54_20,ip_54_21,ip_54_22,ip_54_23,ip_54_24,ip_54_25,ip_54_26,ip_54_27,ip_54_28,ip_54_29,ip_54_30,ip_54_31,ip_54_32,ip_54_33,ip_54_34,ip_54_35,ip_54_36,ip_54_37,ip_54_38,ip_54_39,ip_54_40,ip_54_41,ip_54_42,ip_54_43,ip_54_44,ip_54_45,ip_54_46,ip_54_47,ip_54_48,ip_54_49,ip_54_50,ip_54_51,ip_54_52,ip_54_53,ip_54_54,ip_54_55,ip_54_56,ip_54_57,ip_54_58,ip_54_59,ip_54_60,ip_54_61,ip_54_62,ip_54_63,ip_55_0,ip_55_1,ip_55_2,ip_55_3,ip_55_4,ip_55_5,ip_55_6,ip_55_7,ip_55_8,ip_55_9,ip_55_10,ip_55_11,ip_55_12,ip_55_13,ip_55_14,ip_55_15,ip_55_16,ip_55_17,ip_55_18,ip_55_19,ip_55_20,ip_55_21,ip_55_22,ip_55_23,ip_55_24,ip_55_25,ip_55_26,ip_55_27,ip_55_28,ip_55_29,ip_55_30,ip_55_31,ip_55_32,ip_55_33,ip_55_34,ip_55_35,ip_55_36,ip_55_37,ip_55_38,ip_55_39,ip_55_40,ip_55_41,ip_55_42,ip_55_43,ip_55_44,ip_55_45,ip_55_46,ip_55_47,ip_55_48,ip_55_49,ip_55_50,ip_55_51,ip_55_52,ip_55_53,ip_55_54,ip_55_55,ip_55_56,ip_55_57,ip_55_58,ip_55_59,ip_55_60,ip_55_61,ip_55_62,ip_55_63,ip_56_0,ip_56_1,ip_56_2,ip_56_3,ip_56_4,ip_56_5,ip_56_6,ip_56_7,ip_56_8,ip_56_9,ip_56_10,ip_56_11,ip_56_12,ip_56_13,ip_56_14,ip_56_15,ip_56_16,ip_56_17,ip_56_18,ip_56_19,ip_56_20,ip_56_21,ip_56_22,ip_56_23,ip_56_24,ip_56_25,ip_56_26,ip_56_27,ip_56_28,ip_56_29,ip_56_30,ip_56_31,ip_56_32,ip_56_33,ip_56_34,ip_56_35,ip_56_36,ip_56_37,ip_56_38,ip_56_39,ip_56_40,ip_56_41,ip_56_42,ip_56_43,ip_56_44,ip_56_45,ip_56_46,ip_56_47,ip_56_48,ip_56_49,ip_56_50,ip_56_51,ip_56_52,ip_56_53,ip_56_54,ip_56_55,ip_56_56,ip_56_57,ip_56_58,ip_56_59,ip_56_60,ip_56_61,ip_56_62,ip_56_63,ip_57_0,ip_57_1,ip_57_2,ip_57_3,ip_57_4,ip_57_5,ip_57_6,ip_57_7,ip_57_8,ip_57_9,ip_57_10,ip_57_11,ip_57_12,ip_57_13,ip_57_14,ip_57_15,ip_57_16,ip_57_17,ip_57_18,ip_57_19,ip_57_20,ip_57_21,ip_57_22,ip_57_23,ip_57_24,ip_57_25,ip_57_26,ip_57_27,ip_57_28,ip_57_29,ip_57_30,ip_57_31,ip_57_32,ip_57_33,ip_57_34,ip_57_35,ip_57_36,ip_57_37,ip_57_38,ip_57_39,ip_57_40,ip_57_41,ip_57_42,ip_57_43,ip_57_44,ip_57_45,ip_57_46,ip_57_47,ip_57_48,ip_57_49,ip_57_50,ip_57_51,ip_57_52,ip_57_53,ip_57_54,ip_57_55,ip_57_56,ip_57_57,ip_57_58,ip_57_59,ip_57_60,ip_57_61,ip_57_62,ip_57_63,ip_58_0,ip_58_1,ip_58_2,ip_58_3,ip_58_4,ip_58_5,ip_58_6,ip_58_7,ip_58_8,ip_58_9,ip_58_10,ip_58_11,ip_58_12,ip_58_13,ip_58_14,ip_58_15,ip_58_16,ip_58_17,ip_58_18,ip_58_19,ip_58_20,ip_58_21,ip_58_22,ip_58_23,ip_58_24,ip_58_25,ip_58_26,ip_58_27,ip_58_28,ip_58_29,ip_58_30,ip_58_31,ip_58_32,ip_58_33,ip_58_34,ip_58_35,ip_58_36,ip_58_37,ip_58_38,ip_58_39,ip_58_40,ip_58_41,ip_58_42,ip_58_43,ip_58_44,ip_58_45,ip_58_46,ip_58_47,ip_58_48,ip_58_49,ip_58_50,ip_58_51,ip_58_52,ip_58_53,ip_58_54,ip_58_55,ip_58_56,ip_58_57,ip_58_58,ip_58_59,ip_58_60,ip_58_61,ip_58_62,ip_58_63,ip_59_0,ip_59_1,ip_59_2,ip_59_3,ip_59_4,ip_59_5,ip_59_6,ip_59_7,ip_59_8,ip_59_9,ip_59_10,ip_59_11,ip_59_12,ip_59_13,ip_59_14,ip_59_15,ip_59_16,ip_59_17,ip_59_18,ip_59_19,ip_59_20,ip_59_21,ip_59_22,ip_59_23,ip_59_24,ip_59_25,ip_59_26,ip_59_27,ip_59_28,ip_59_29,ip_59_30,ip_59_31,ip_59_32,ip_59_33,ip_59_34,ip_59_35,ip_59_36,ip_59_37,ip_59_38,ip_59_39,ip_59_40,ip_59_41,ip_59_42,ip_59_43,ip_59_44,ip_59_45,ip_59_46,ip_59_47,ip_59_48,ip_59_49,ip_59_50,ip_59_51,ip_59_52,ip_59_53,ip_59_54,ip_59_55,ip_59_56,ip_59_57,ip_59_58,ip_59_59,ip_59_60,ip_59_61,ip_59_62,ip_59_63,ip_60_0,ip_60_1,ip_60_2,ip_60_3,ip_60_4,ip_60_5,ip_60_6,ip_60_7,ip_60_8,ip_60_9,ip_60_10,ip_60_11,ip_60_12,ip_60_13,ip_60_14,ip_60_15,ip_60_16,ip_60_17,ip_60_18,ip_60_19,ip_60_20,ip_60_21,ip_60_22,ip_60_23,ip_60_24,ip_60_25,ip_60_26,ip_60_27,ip_60_28,ip_60_29,ip_60_30,ip_60_31,ip_60_32,ip_60_33,ip_60_34,ip_60_35,ip_60_36,ip_60_37,ip_60_38,ip_60_39,ip_60_40,ip_60_41,ip_60_42,ip_60_43,ip_60_44,ip_60_45,ip_60_46,ip_60_47,ip_60_48,ip_60_49,ip_60_50,ip_60_51,ip_60_52,ip_60_53,ip_60_54,ip_60_55,ip_60_56,ip_60_57,ip_60_58,ip_60_59,ip_60_60,ip_60_61,ip_60_62,ip_60_63,ip_61_0,ip_61_1,ip_61_2,ip_61_3,ip_61_4,ip_61_5,ip_61_6,ip_61_7,ip_61_8,ip_61_9,ip_61_10,ip_61_11,ip_61_12,ip_61_13,ip_61_14,ip_61_15,ip_61_16,ip_61_17,ip_61_18,ip_61_19,ip_61_20,ip_61_21,ip_61_22,ip_61_23,ip_61_24,ip_61_25,ip_61_26,ip_61_27,ip_61_28,ip_61_29,ip_61_30,ip_61_31,ip_61_32,ip_61_33,ip_61_34,ip_61_35,ip_61_36,ip_61_37,ip_61_38,ip_61_39,ip_61_40,ip_61_41,ip_61_42,ip_61_43,ip_61_44,ip_61_45,ip_61_46,ip_61_47,ip_61_48,ip_61_49,ip_61_50,ip_61_51,ip_61_52,ip_61_53,ip_61_54,ip_61_55,ip_61_56,ip_61_57,ip_61_58,ip_61_59,ip_61_60,ip_61_61,ip_61_62,ip_61_63,ip_62_0,ip_62_1,ip_62_2,ip_62_3,ip_62_4,ip_62_5,ip_62_6,ip_62_7,ip_62_8,ip_62_9,ip_62_10,ip_62_11,ip_62_12,ip_62_13,ip_62_14,ip_62_15,ip_62_16,ip_62_17,ip_62_18,ip_62_19,ip_62_20,ip_62_21,ip_62_22,ip_62_23,ip_62_24,ip_62_25,ip_62_26,ip_62_27,ip_62_28,ip_62_29,ip_62_30,ip_62_31,ip_62_32,ip_62_33,ip_62_34,ip_62_35,ip_62_36,ip_62_37,ip_62_38,ip_62_39,ip_62_40,ip_62_41,ip_62_42,ip_62_43,ip_62_44,ip_62_45,ip_62_46,ip_62_47,ip_62_48,ip_62_49,ip_62_50,ip_62_51,ip_62_52,ip_62_53,ip_62_54,ip_62_55,ip_62_56,ip_62_57,ip_62_58,ip_62_59,ip_62_60,ip_62_61,ip_62_62,ip_62_63,ip_63_0,ip_63_1,ip_63_2,ip_63_3,ip_63_4,ip_63_5,ip_63_6,ip_63_7,ip_63_8,ip_63_9,ip_63_10,ip_63_11,ip_63_12,ip_63_13,ip_63_14,ip_63_15,ip_63_16,ip_63_17,ip_63_18,ip_63_19,ip_63_20,ip_63_21,ip_63_22,ip_63_23,ip_63_24,ip_63_25,ip_63_26,ip_63_27,ip_63_28,ip_63_29,ip_63_30,ip_63_31,ip_63_32,ip_63_33,ip_63_34,ip_63_35,ip_63_36,ip_63_37,ip_63_38,ip_63_39,ip_63_40,ip_63_41,ip_63_42,ip_63_43,ip_63_44,ip_63_45,ip_63_46,ip_63_47,ip_63_48,ip_63_49,ip_63_50,ip_63_51,ip_63_52,ip_63_53,ip_63_54,ip_63_55,ip_63_56,ip_63_57,ip_63_58,ip_63_59,ip_63_60,ip_63_61,ip_63_62,ip_63_63;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117,p118,p119,p120,p121,p122,p123,p124,p125,p126,p127,p128,p129,p130,p131,p132,p133,p134,p135,p136,p137,p138,p139,p140,p141,p142,p143,p144,p145,p146,p147,p148,p149,p150,p151,p152,p153,p154,p155,p156,p157,p158,p159,p160,p161,p162,p163,p164,p165,p166,p167,p168,p169,p170,p171,p172,p173,p174,p175,p176,p177,p178,p179,p180,p181,p182,p183,p184,p185,p186,p187,p188,p189,p190,p191,p192,p193,p194,p195,p196,p197,p198,p199,p200,p201,p202,p203,p204,p205,p206,p207,p208,p209,p210,p211,p212,p213,p214,p215,p216,p217,p218,p219,p220,p221,p222,p223,p224,p225,p226,p227,p228,p229,p230,p231,p232,p233,p234,p235,p236,p237,p238,p239,p240,p241,p242,p243,p244,p245,p246,p247,p248,p249,p250,p251,p252,p253,p254,p255,p256,p257,p258,p259,p260,p261,p262,p263,p264,p265,p266,p267,p268,p269,p270,p271,p272,p273,p274,p275,p276,p277,p278,p279,p280,p281,p282,p283,p284,p285,p286,p287,p288,p289,p290,p291,p292,p293,p294,p295,p296,p297,p298,p299,p300,p301,p302,p303,p304,p305,p306,p307,p308,p309,p310,p311,p312,p313,p314,p315,p316,p317,p318,p319,p320,p321,p322,p323,p324,p325,p326,p327,p328,p329,p330,p331,p332,p333,p334,p335,p336,p337,p338,p339,p340,p341,p342,p343,p344,p345,p346,p347,p348,p349,p350,p351,p352,p353,p354,p355,p356,p357,p358,p359,p360,p361,p362,p363,p364,p365,p366,p367,p368,p369,p370,p371,p372,p373,p374,p375,p376,p377,p378,p379,p380,p381,p382,p383,p384,p385,p386,p387,p388,p389,p390,p391,p392,p393,p394,p395,p396,p397,p398,p399,p400,p401,p402,p403,p404,p405,p406,p407,p408,p409,p410,p411,p412,p413,p414,p415,p416,p417,p418,p419,p420,p421,p422,p423,p424,p425,p426,p427,p428,p429,p430,p431,p432,p433,p434,p435,p436,p437,p438,p439,p440,p441,p442,p443,p444,p445,p446,p447,p448,p449,p450,p451,p452,p453,p454,p455,p456,p457,p458,p459,p460,p461,p462,p463,p464,p465,p466,p467,p468,p469,p470,p471,p472,p473,p474,p475,p476,p477,p478,p479,p480,p481,p482,p483,p484,p485,p486,p487,p488,p489,p490,p491,p492,p493,p494,p495,p496,p497,p498,p499,p500,p501,p502,p503,p504,p505,p506,p507,p508,p509,p510,p511,p512,p513,p514,p515,p516,p517,p518,p519,p520,p521,p522,p523,p524,p525,p526,p527,p528,p529,p530,p531,p532,p533,p534,p535,p536,p537,p538,p539,p540,p541,p542,p543,p544,p545,p546,p547,p548,p549,p550,p551,p552,p553,p554,p555,p556,p557,p558,p559,p560,p561,p562,p563,p564,p565,p566,p567,p568,p569,p570,p571,p572,p573,p574,p575,p576,p577,p578,p579,p580,p581,p582,p583,p584,p585,p586,p587,p588,p589,p590,p591,p592,p593,p594,p595,p596,p597,p598,p599,p600,p601,p602,p603,p604,p605,p606,p607,p608,p609,p610,p611,p612,p613,p614,p615,p616,p617,p618,p619,p620,p621,p622,p623,p624,p625,p626,p627,p628,p629,p630,p631,p632,p633,p634,p635,p636,p637,p638,p639,p640,p641,p642,p643,p644,p645,p646,p647,p648,p649,p650,p651,p652,p653,p654,p655,p656,p657,p658,p659,p660,p661,p662,p663,p664,p665,p666,p667,p668,p669,p670,p671,p672,p673,p674,p675,p676,p677,p678,p679,p680,p681,p682,p683,p684,p685,p686,p687,p688,p689,p690,p691,p692,p693,p694,p695,p696,p697,p698,p699,p700,p701,p702,p703,p704,p705,p706,p707,p708,p709,p710,p711,p712,p713,p714,p715,p716,p717,p718,p719,p720,p721,p722,p723,p724,p725,p726,p727,p728,p729,p730,p731,p732,p733,p734,p735,p736,p737,p738,p739,p740,p741,p742,p743,p744,p745,p746,p747,p748,p749,p750,p751,p752,p753,p754,p755,p756,p757,p758,p759,p760,p761,p762,p763,p764,p765,p766,p767,p768,p769,p770,p771,p772,p773,p774,p775,p776,p777,p778,p779,p780,p781,p782,p783,p784,p785,p786,p787,p788,p789,p790,p791,p792,p793,p794,p795,p796,p797,p798,p799,p800,p801,p802,p803,p804,p805,p806,p807,p808,p809,p810,p811,p812,p813,p814,p815,p816,p817,p818,p819,p820,p821,p822,p823,p824,p825,p826,p827,p828,p829,p830,p831,p832,p833,p834,p835,p836,p837,p838,p839,p840,p841,p842,p843,p844,p845,p846,p847,p848,p849,p850,p851,p852,p853,p854,p855,p856,p857,p858,p859,p860,p861,p862,p863,p864,p865,p866,p867,p868,p869,p870,p871,p872,p873,p874,p875,p876,p877,p878,p879,p880,p881,p882,p883,p884,p885,p886,p887,p888,p889,p890,p891,p892,p893,p894,p895,p896,p897,p898,p899,p900,p901,p902,p903,p904,p905,p906,p907,p908,p909,p910,p911,p912,p913,p914,p915,p916,p917,p918,p919,p920,p921,p922,p923,p924,p925,p926,p927,p928,p929,p930,p931,p932,p933,p934,p935,p936,p937,p938,p939,p940,p941,p942,p943,p944,p945,p946,p947,p948,p949,p950,p951,p952,p953,p954,p955,p956,p957,p958,p959,p960,p961,p962,p963,p964,p965,p966,p967,p968,p969,p970,p971,p972,p973,p974,p975,p976,p977,p978,p979,p980,p981,p982,p983,p984,p985,p986,p987,p988,p989,p990,p991,p992,p993,p994,p995,p996,p997,p998,p999,p1000,p1001,p1002,p1003,p1004,p1005,p1006,p1007,p1008,p1009,p1010,p1011,p1012,p1013,p1014,p1015,p1016,p1017,p1018,p1019,p1020,p1021,p1022,p1023,p1024,p1025,p1026,p1027,p1028,p1029,p1030,p1031,p1032,p1033,p1034,p1035,p1036,p1037,p1038,p1039,p1040,p1041,p1042,p1043,p1044,p1045,p1046,p1047,p1048,p1049,p1050,p1051,p1052,p1053,p1054,p1055,p1056,p1057,p1058,p1059,p1060,p1061,p1062,p1063,p1064,p1065,p1066,p1067,p1068,p1069,p1070,p1071,p1072,p1073,p1074,p1075,p1076,p1077,p1078,p1079,p1080,p1081,p1082,p1083,p1084,p1085,p1086,p1087,p1088,p1089,p1090,p1091,p1092,p1093,p1094,p1095,p1096,p1097,p1098,p1099,p1100,p1101,p1102,p1103,p1104,p1105,p1106,p1107,p1108,p1109,p1110,p1111,p1112,p1113,p1114,p1115,p1116,p1117,p1118,p1119,p1120,p1121,p1122,p1123,p1124,p1125,p1126,p1127,p1128,p1129,p1130,p1131,p1132,p1133,p1134,p1135,p1136,p1137,p1138,p1139,p1140,p1141,p1142,p1143,p1144,p1145,p1146,p1147,p1148,p1149,p1150,p1151,p1152,p1153,p1154,p1155,p1156,p1157,p1158,p1159,p1160,p1161,p1162,p1163,p1164,p1165,p1166,p1167,p1168,p1169,p1170,p1171,p1172,p1173,p1174,p1175,p1176,p1177,p1178,p1179,p1180,p1181,p1182,p1183,p1184,p1185,p1186,p1187,p1188,p1189,p1190,p1191,p1192,p1193,p1194,p1195,p1196,p1197,p1198,p1199,p1200,p1201,p1202,p1203,p1204,p1205,p1206,p1207,p1208,p1209,p1210,p1211,p1212,p1213,p1214,p1215,p1216,p1217,p1218,p1219,p1220,p1221,p1222,p1223,p1224,p1225,p1226,p1227,p1228,p1229,p1230,p1231,p1232,p1233,p1234,p1235,p1236,p1237,p1238,p1239,p1240,p1241,p1242,p1243,p1244,p1245,p1246,p1247,p1248,p1249,p1250,p1251,p1252,p1253,p1254,p1255,p1256,p1257,p1258,p1259,p1260,p1261,p1262,p1263,p1264,p1265,p1266,p1267,p1268,p1269,p1270,p1271,p1272,p1273,p1274,p1275,p1276,p1277,p1278,p1279,p1280,p1281,p1282,p1283,p1284,p1285,p1286,p1287,p1288,p1289,p1290,p1291,p1292,p1293,p1294,p1295,p1296,p1297,p1298,p1299,p1300,p1301,p1302,p1303,p1304,p1305,p1306,p1307,p1308,p1309,p1310,p1311,p1312,p1313,p1314,p1315,p1316,p1317,p1318,p1319,p1320,p1321,p1322,p1323,p1324,p1325,p1326,p1327,p1328,p1329,p1330,p1331,p1332,p1333,p1334,p1335,p1336,p1337,p1338,p1339,p1340,p1341,p1342,p1343,p1344,p1345,p1346,p1347,p1348,p1349,p1350,p1351,p1352,p1353,p1354,p1355,p1356,p1357,p1358,p1359,p1360,p1361,p1362,p1363,p1364,p1365,p1366,p1367,p1368,p1369,p1370,p1371,p1372,p1373,p1374,p1375,p1376,p1377,p1378,p1379,p1380,p1381,p1382,p1383,p1384,p1385,p1386,p1387,p1388,p1389,p1390,p1391,p1392,p1393,p1394,p1395,p1396,p1397,p1398,p1399,p1400,p1401,p1402,p1403,p1404,p1405,p1406,p1407,p1408,p1409,p1410,p1411,p1412,p1413,p1414,p1415,p1416,p1417,p1418,p1419,p1420,p1421,p1422,p1423,p1424,p1425,p1426,p1427,p1428,p1429,p1430,p1431,p1432,p1433,p1434,p1435,p1436,p1437,p1438,p1439,p1440,p1441,p1442,p1443,p1444,p1445,p1446,p1447,p1448,p1449,p1450,p1451,p1452,p1453,p1454,p1455,p1456,p1457,p1458,p1459,p1460,p1461,p1462,p1463,p1464,p1465,p1466,p1467,p1468,p1469,p1470,p1471,p1472,p1473,p1474,p1475,p1476,p1477,p1478,p1479,p1480,p1481,p1482,p1483,p1484,p1485,p1486,p1487,p1488,p1489,p1490,p1491,p1492,p1493,p1494,p1495,p1496,p1497,p1498,p1499,p1500,p1501,p1502,p1503,p1504,p1505,p1506,p1507,p1508,p1509,p1510,p1511,p1512,p1513,p1514,p1515,p1516,p1517,p1518,p1519,p1520,p1521,p1522,p1523,p1524,p1525,p1526,p1527,p1528,p1529,p1530,p1531,p1532,p1533,p1534,p1535,p1536,p1537,p1538,p1539,p1540,p1541,p1542,p1543,p1544,p1545,p1546,p1547,p1548,p1549,p1550,p1551,p1552,p1553,p1554,p1555,p1556,p1557,p1558,p1559,p1560,p1561,p1562,p1563,p1564,p1565,p1566,p1567,p1568,p1569,p1570,p1571,p1572,p1573,p1574,p1575,p1576,p1577,p1578,p1579,p1580,p1581,p1582,p1583,p1584,p1585,p1586,p1587,p1588,p1589,p1590,p1591,p1592,p1593,p1594,p1595,p1596,p1597,p1598,p1599,p1600,p1601,p1602,p1603,p1604,p1605,p1606,p1607,p1608,p1609,p1610,p1611,p1612,p1613,p1614,p1615,p1616,p1617,p1618,p1619,p1620,p1621,p1622,p1623,p1624,p1625,p1626,p1627,p1628,p1629,p1630,p1631,p1632,p1633,p1634,p1635,p1636,p1637,p1638,p1639,p1640,p1641,p1642,p1643,p1644,p1645,p1646,p1647,p1648,p1649,p1650,p1651,p1652,p1653,p1654,p1655,p1656,p1657,p1658,p1659,p1660,p1661,p1662,p1663,p1664,p1665,p1666,p1667,p1668,p1669,p1670,p1671,p1672,p1673,p1674,p1675,p1676,p1677,p1678,p1679,p1680,p1681,p1682,p1683,p1684,p1685,p1686,p1687,p1688,p1689,p1690,p1691,p1692,p1693,p1694,p1695,p1696,p1697,p1698,p1699,p1700,p1701,p1702,p1703,p1704,p1705,p1706,p1707,p1708,p1709,p1710,p1711,p1712,p1713,p1714,p1715,p1716,p1717,p1718,p1719,p1720,p1721,p1722,p1723,p1724,p1725,p1726,p1727,p1728,p1729,p1730,p1731,p1732,p1733,p1734,p1735,p1736,p1737,p1738,p1739,p1740,p1741,p1742,p1743,p1744,p1745,p1746,p1747,p1748,p1749,p1750,p1751,p1752,p1753,p1754,p1755,p1756,p1757,p1758,p1759,p1760,p1761,p1762,p1763,p1764,p1765,p1766,p1767,p1768,p1769,p1770,p1771,p1772,p1773,p1774,p1775,p1776,p1777,p1778,p1779,p1780,p1781,p1782,p1783,p1784,p1785,p1786,p1787,p1788,p1789,p1790,p1791,p1792,p1793,p1794,p1795,p1796,p1797,p1798,p1799,p1800,p1801,p1802,p1803,p1804,p1805,p1806,p1807,p1808,p1809,p1810,p1811,p1812,p1813,p1814,p1815,p1816,p1817,p1818,p1819,p1820,p1821,p1822,p1823,p1824,p1825,p1826,p1827,p1828,p1829,p1830,p1831,p1832,p1833,p1834,p1835,p1836,p1837,p1838,p1839,p1840,p1841,p1842,p1843,p1844,p1845,p1846,p1847,p1848,p1849,p1850,p1851,p1852,p1853,p1854,p1855,p1856,p1857,p1858,p1859,p1860,p1861,p1862,p1863,p1864,p1865,p1866,p1867,p1868,p1869,p1870,p1871,p1872,p1873,p1874,p1875,p1876,p1877,p1878,p1879,p1880,p1881,p1882,p1883,p1884,p1885,p1886,p1887,p1888,p1889,p1890,p1891,p1892,p1893,p1894,p1895,p1896,p1897,p1898,p1899,p1900,p1901,p1902,p1903,p1904,p1905,p1906,p1907,p1908,p1909,p1910,p1911,p1912,p1913,p1914,p1915,p1916,p1917,p1918,p1919,p1920,p1921,p1922,p1923,p1924,p1925,p1926,p1927,p1928,p1929,p1930,p1931,p1932,p1933,p1934,p1935,p1936,p1937,p1938,p1939,p1940,p1941,p1942,p1943,p1944,p1945,p1946,p1947,p1948,p1949,p1950,p1951,p1952,p1953,p1954,p1955,p1956,p1957,p1958,p1959,p1960,p1961,p1962,p1963,p1964,p1965,p1966,p1967,p1968,p1969,p1970,p1971,p1972,p1973,p1974,p1975,p1976,p1977,p1978,p1979,p1980,p1981,p1982,p1983,p1984,p1985,p1986,p1987,p1988,p1989,p1990,p1991,p1992,p1993,p1994,p1995,p1996,p1997,p1998,p1999,p2000,p2001,p2002,p2003,p2004,p2005,p2006,p2007,p2008,p2009,p2010,p2011,p2012,p2013,p2014,p2015,p2016,p2017,p2018,p2019,p2020,p2021,p2022,p2023,p2024,p2025,p2026,p2027,p2028,p2029,p2030,p2031,p2032,p2033,p2034,p2035,p2036,p2037,p2038,p2039,p2040,p2041,p2042,p2043,p2044,p2045,p2046,p2047,p2048,p2049,p2050,p2051,p2052,p2053,p2054,p2055,p2056,p2057,p2058,p2059,p2060,p2061,p2062,p2063,p2064,p2065,p2066,p2067,p2068,p2069,p2070,p2071,p2072,p2073,p2074,p2075,p2076,p2077,p2078,p2079,p2080,p2081,p2082,p2083,p2084,p2085,p2086,p2087,p2088,p2089,p2090,p2091,p2092,p2093,p2094,p2095,p2096,p2097,p2098,p2099,p2100,p2101,p2102,p2103,p2104,p2105,p2106,p2107,p2108,p2109,p2110,p2111,p2112,p2113,p2114,p2115,p2116,p2117,p2118,p2119,p2120,p2121,p2122,p2123,p2124,p2125,p2126,p2127,p2128,p2129,p2130,p2131,p2132,p2133,p2134,p2135,p2136,p2137,p2138,p2139,p2140,p2141,p2142,p2143,p2144,p2145,p2146,p2147,p2148,p2149,p2150,p2151,p2152,p2153,p2154,p2155,p2156,p2157,p2158,p2159,p2160,p2161,p2162,p2163,p2164,p2165,p2166,p2167,p2168,p2169,p2170,p2171,p2172,p2173,p2174,p2175,p2176,p2177,p2178,p2179,p2180,p2181,p2182,p2183,p2184,p2185,p2186,p2187,p2188,p2189,p2190,p2191,p2192,p2193,p2194,p2195,p2196,p2197,p2198,p2199,p2200,p2201,p2202,p2203,p2204,p2205,p2206,p2207,p2208,p2209,p2210,p2211,p2212,p2213,p2214,p2215,p2216,p2217,p2218,p2219,p2220,p2221,p2222,p2223,p2224,p2225,p2226,p2227,p2228,p2229,p2230,p2231,p2232,p2233,p2234,p2235,p2236,p2237,p2238,p2239,p2240,p2241,p2242,p2243,p2244,p2245,p2246,p2247,p2248,p2249,p2250,p2251,p2252,p2253,p2254,p2255,p2256,p2257,p2258,p2259,p2260,p2261,p2262,p2263,p2264,p2265,p2266,p2267,p2268,p2269,p2270,p2271,p2272,p2273,p2274,p2275,p2276,p2277,p2278,p2279,p2280,p2281,p2282,p2283,p2284,p2285,p2286,p2287,p2288,p2289,p2290,p2291,p2292,p2293,p2294,p2295,p2296,p2297,p2298,p2299,p2300,p2301,p2302,p2303,p2304,p2305,p2306,p2307,p2308,p2309,p2310,p2311,p2312,p2313,p2314,p2315,p2316,p2317,p2318,p2319,p2320,p2321,p2322,p2323,p2324,p2325,p2326,p2327,p2328,p2329,p2330,p2331,p2332,p2333,p2334,p2335,p2336,p2337,p2338,p2339,p2340,p2341,p2342,p2343,p2344,p2345,p2346,p2347,p2348,p2349,p2350,p2351,p2352,p2353,p2354,p2355,p2356,p2357,p2358,p2359,p2360,p2361,p2362,p2363,p2364,p2365,p2366,p2367,p2368,p2369,p2370,p2371,p2372,p2373,p2374,p2375,p2376,p2377,p2378,p2379,p2380,p2381,p2382,p2383,p2384,p2385,p2386,p2387,p2388,p2389,p2390,p2391,p2392,p2393,p2394,p2395,p2396,p2397,p2398,p2399,p2400,p2401,p2402,p2403,p2404,p2405,p2406,p2407,p2408,p2409,p2410,p2411,p2412,p2413,p2414,p2415,p2416,p2417,p2418,p2419,p2420,p2421,p2422,p2423,p2424,p2425,p2426,p2427,p2428,p2429,p2430,p2431,p2432,p2433,p2434,p2435,p2436,p2437,p2438,p2439,p2440,p2441,p2442,p2443,p2444,p2445,p2446,p2447,p2448,p2449,p2450,p2451,p2452,p2453,p2454,p2455,p2456,p2457,p2458,p2459,p2460,p2461,p2462,p2463,p2464,p2465,p2466,p2467,p2468,p2469,p2470,p2471,p2472,p2473,p2474,p2475,p2476,p2477,p2478,p2479,p2480,p2481,p2482,p2483,p2484,p2485,p2486,p2487,p2488,p2489,p2490,p2491,p2492,p2493,p2494,p2495,p2496,p2497,p2498,p2499,p2500,p2501,p2502,p2503,p2504,p2505,p2506,p2507,p2508,p2509,p2510,p2511,p2512,p2513,p2514,p2515,p2516,p2517,p2518,p2519,p2520,p2521,p2522,p2523,p2524,p2525,p2526,p2527,p2528,p2529,p2530,p2531,p2532,p2533,p2534,p2535,p2536,p2537,p2538,p2539,p2540,p2541,p2542,p2543,p2544,p2545,p2546,p2547,p2548,p2549,p2550,p2551,p2552,p2553,p2554,p2555,p2556,p2557,p2558,p2559,p2560,p2561,p2562,p2563,p2564,p2565,p2566,p2567,p2568,p2569,p2570,p2571,p2572,p2573,p2574,p2575,p2576,p2577,p2578,p2579,p2580,p2581,p2582,p2583,p2584,p2585,p2586,p2587,p2588,p2589,p2590,p2591,p2592,p2593,p2594,p2595,p2596,p2597,p2598,p2599,p2600,p2601,p2602,p2603,p2604,p2605,p2606,p2607,p2608,p2609,p2610,p2611,p2612,p2613,p2614,p2615,p2616,p2617,p2618,p2619,p2620,p2621,p2622,p2623,p2624,p2625,p2626,p2627,p2628,p2629,p2630,p2631,p2632,p2633,p2634,p2635,p2636,p2637,p2638,p2639,p2640,p2641,p2642,p2643,p2644,p2645,p2646,p2647,p2648,p2649,p2650,p2651,p2652,p2653,p2654,p2655,p2656,p2657,p2658,p2659,p2660,p2661,p2662,p2663,p2664,p2665,p2666,p2667,p2668,p2669,p2670,p2671,p2672,p2673,p2674,p2675,p2676,p2677,p2678,p2679,p2680,p2681,p2682,p2683,p2684,p2685,p2686,p2687,p2688,p2689,p2690,p2691,p2692,p2693,p2694,p2695,p2696,p2697,p2698,p2699,p2700,p2701,p2702,p2703,p2704,p2705,p2706,p2707,p2708,p2709,p2710,p2711,p2712,p2713,p2714,p2715,p2716,p2717,p2718,p2719,p2720,p2721,p2722,p2723,p2724,p2725,p2726,p2727,p2728,p2729,p2730,p2731,p2732,p2733,p2734,p2735,p2736,p2737,p2738,p2739,p2740,p2741,p2742,p2743,p2744,p2745,p2746,p2747,p2748,p2749,p2750,p2751,p2752,p2753,p2754,p2755,p2756,p2757,p2758,p2759,p2760,p2761,p2762,p2763,p2764,p2765,p2766,p2767,p2768,p2769,p2770,p2771,p2772,p2773,p2774,p2775,p2776,p2777,p2778,p2779,p2780,p2781,p2782,p2783,p2784,p2785,p2786,p2787,p2788,p2789,p2790,p2791,p2792,p2793,p2794,p2795,p2796,p2797,p2798,p2799,p2800,p2801,p2802,p2803,p2804,p2805,p2806,p2807,p2808,p2809,p2810,p2811,p2812,p2813,p2814,p2815,p2816,p2817,p2818,p2819,p2820,p2821,p2822,p2823,p2824,p2825,p2826,p2827,p2828,p2829,p2830,p2831,p2832,p2833,p2834,p2835,p2836,p2837,p2838,p2839,p2840,p2841,p2842,p2843,p2844,p2845,p2846,p2847,p2848,p2849,p2850,p2851,p2852,p2853,p2854,p2855,p2856,p2857,p2858,p2859,p2860,p2861,p2862,p2863,p2864,p2865,p2866,p2867,p2868,p2869,p2870,p2871,p2872,p2873,p2874,p2875,p2876,p2877,p2878,p2879,p2880,p2881,p2882,p2883,p2884,p2885,p2886,p2887,p2888,p2889,p2890,p2891,p2892,p2893,p2894,p2895,p2896,p2897,p2898,p2899,p2900,p2901,p2902,p2903,p2904,p2905,p2906,p2907,p2908,p2909,p2910,p2911,p2912,p2913,p2914,p2915,p2916,p2917,p2918,p2919,p2920,p2921,p2922,p2923,p2924,p2925,p2926,p2927,p2928,p2929,p2930,p2931,p2932,p2933,p2934,p2935,p2936,p2937,p2938,p2939,p2940,p2941,p2942,p2943,p2944,p2945,p2946,p2947,p2948,p2949,p2950,p2951,p2952,p2953,p2954,p2955,p2956,p2957,p2958,p2959,p2960,p2961,p2962,p2963,p2964,p2965,p2966,p2967,p2968,p2969,p2970,p2971,p2972,p2973,p2974,p2975,p2976,p2977,p2978,p2979,p2980,p2981,p2982,p2983,p2984,p2985,p2986,p2987,p2988,p2989,p2990,p2991,p2992,p2993,p2994,p2995,p2996,p2997,p2998,p2999,p3000,p3001,p3002,p3003,p3004,p3005,p3006,p3007,p3008,p3009,p3010,p3011,p3012,p3013,p3014,p3015,p3016,p3017,p3018,p3019,p3020,p3021,p3022,p3023,p3024,p3025,p3026,p3027,p3028,p3029,p3030,p3031,p3032,p3033,p3034,p3035,p3036,p3037,p3038,p3039,p3040,p3041,p3042,p3043,p3044,p3045,p3046,p3047,p3048,p3049,p3050,p3051,p3052,p3053,p3054,p3055,p3056,p3057,p3058,p3059,p3060,p3061,p3062,p3063,p3064,p3065,p3066,p3067,p3068,p3069,p3070,p3071,p3072,p3073,p3074,p3075,p3076,p3077,p3078,p3079,p3080,p3081,p3082,p3083,p3084,p3085,p3086,p3087,p3088,p3089,p3090,p3091,p3092,p3093,p3094,p3095,p3096,p3097,p3098,p3099,p3100,p3101,p3102,p3103,p3104,p3105,p3106,p3107,p3108,p3109,p3110,p3111,p3112,p3113,p3114,p3115,p3116,p3117,p3118,p3119,p3120,p3121,p3122,p3123,p3124,p3125,p3126,p3127,p3128,p3129,p3130,p3131,p3132,p3133,p3134,p3135,p3136,p3137,p3138,p3139,p3140,p3141,p3142,p3143,p3144,p3145,p3146,p3147,p3148,p3149,p3150,p3151,p3152,p3153,p3154,p3155,p3156,p3157,p3158,p3159,p3160,p3161,p3162,p3163,p3164,p3165,p3166,p3167,p3168,p3169,p3170,p3171,p3172,p3173,p3174,p3175,p3176,p3177,p3178,p3179,p3180,p3181,p3182,p3183,p3184,p3185,p3186,p3187,p3188,p3189,p3190,p3191,p3192,p3193,p3194,p3195,p3196,p3197,p3198,p3199,p3200,p3201,p3202,p3203,p3204,p3205,p3206,p3207,p3208,p3209,p3210,p3211,p3212,p3213,p3214,p3215,p3216,p3217,p3218,p3219,p3220,p3221,p3222,p3223,p3224,p3225,p3226,p3227,p3228,p3229,p3230,p3231,p3232,p3233,p3234,p3235,p3236,p3237,p3238,p3239,p3240,p3241,p3242,p3243,p3244,p3245,p3246,p3247,p3248,p3249,p3250,p3251,p3252,p3253,p3254,p3255,p3256,p3257,p3258,p3259,p3260,p3261,p3262,p3263,p3264,p3265,p3266,p3267,p3268,p3269,p3270,p3271,p3272,p3273,p3274,p3275,p3276,p3277,p3278,p3279,p3280,p3281,p3282,p3283,p3284,p3285,p3286,p3287,p3288,p3289,p3290,p3291,p3292,p3293,p3294,p3295,p3296,p3297,p3298,p3299,p3300,p3301,p3302,p3303,p3304,p3305,p3306,p3307,p3308,p3309,p3310,p3311,p3312,p3313,p3314,p3315,p3316,p3317,p3318,p3319,p3320,p3321,p3322,p3323,p3324,p3325,p3326,p3327,p3328,p3329,p3330,p3331,p3332,p3333,p3334,p3335,p3336,p3337,p3338,p3339,p3340,p3341,p3342,p3343,p3344,p3345,p3346,p3347,p3348,p3349,p3350,p3351,p3352,p3353,p3354,p3355,p3356,p3357,p3358,p3359,p3360,p3361,p3362,p3363,p3364,p3365,p3366,p3367,p3368,p3369,p3370,p3371,p3372,p3373,p3374,p3375,p3376,p3377,p3378,p3379,p3380,p3381,p3382,p3383,p3384,p3385,p3386,p3387,p3388,p3389,p3390,p3391,p3392,p3393,p3394,p3395,p3396,p3397,p3398,p3399,p3400,p3401,p3402,p3403,p3404,p3405,p3406,p3407,p3408,p3409,p3410,p3411,p3412,p3413,p3414,p3415,p3416,p3417,p3418,p3419,p3420,p3421,p3422,p3423,p3424,p3425,p3426,p3427,p3428,p3429,p3430,p3431,p3432,p3433,p3434,p3435,p3436,p3437,p3438,p3439,p3440,p3441,p3442,p3443,p3444,p3445,p3446,p3447,p3448,p3449,p3450,p3451,p3452,p3453,p3454,p3455,p3456,p3457,p3458,p3459,p3460,p3461,p3462,p3463,p3464,p3465,p3466,p3467,p3468,p3469,p3470,p3471,p3472,p3473,p3474,p3475,p3476,p3477,p3478,p3479,p3480,p3481,p3482,p3483,p3484,p3485,p3486,p3487,p3488,p3489,p3490,p3491,p3492,p3493,p3494,p3495,p3496,p3497,p3498,p3499,p3500,p3501,p3502,p3503,p3504,p3505,p3506,p3507,p3508,p3509,p3510,p3511,p3512,p3513,p3514,p3515,p3516,p3517,p3518,p3519,p3520,p3521,p3522,p3523,p3524,p3525,p3526,p3527,p3528,p3529,p3530,p3531,p3532,p3533,p3534,p3535,p3536,p3537,p3538,p3539,p3540,p3541,p3542,p3543,p3544,p3545,p3546,p3547,p3548,p3549,p3550,p3551,p3552,p3553,p3554,p3555,p3556,p3557,p3558,p3559,p3560,p3561,p3562,p3563,p3564,p3565,p3566,p3567,p3568,p3569,p3570,p3571,p3572,p3573,p3574,p3575,p3576,p3577,p3578,p3579,p3580,p3581,p3582,p3583,p3584,p3585,p3586,p3587,p3588,p3589,p3590,p3591,p3592,p3593,p3594,p3595,p3596,p3597,p3598,p3599,p3600,p3601,p3602,p3603,p3604,p3605,p3606,p3607,p3608,p3609,p3610,p3611,p3612,p3613,p3614,p3615,p3616,p3617,p3618,p3619,p3620,p3621,p3622,p3623,p3624,p3625,p3626,p3627,p3628,p3629,p3630,p3631,p3632,p3633,p3634,p3635,p3636,p3637,p3638,p3639,p3640,p3641,p3642,p3643,p3644,p3645,p3646,p3647,p3648,p3649,p3650,p3651,p3652,p3653,p3654,p3655,p3656,p3657,p3658,p3659,p3660,p3661,p3662,p3663,p3664,p3665,p3666,p3667,p3668,p3669,p3670,p3671,p3672,p3673,p3674,p3675,p3676,p3677,p3678,p3679,p3680,p3681,p3682,p3683,p3684,p3685,p3686,p3687,p3688,p3689,p3690,p3691,p3692,p3693,p3694,p3695,p3696,p3697,p3698,p3699,p3700,p3701,p3702,p3703,p3704,p3705,p3706,p3707,p3708,p3709,p3710,p3711,p3712,p3713,p3714,p3715,p3716,p3717,p3718,p3719,p3720,p3721,p3722,p3723,p3724,p3725,p3726,p3727,p3728,p3729,p3730,p3731,p3732,p3733,p3734,p3735,p3736,p3737,p3738,p3739,p3740,p3741,p3742,p3743,p3744,p3745,p3746,p3747,p3748,p3749,p3750,p3751,p3752,p3753,p3754,p3755,p3756,p3757,p3758,p3759,p3760,p3761,p3762,p3763,p3764,p3765,p3766,p3767,p3768,p3769,p3770,p3771,p3772,p3773,p3774,p3775,p3776,p3777,p3778,p3779,p3780,p3781,p3782,p3783,p3784,p3785,p3786,p3787,p3788,p3789,p3790,p3791,p3792,p3793,p3794,p3795,p3796,p3797,p3798,p3799,p3800,p3801,p3802,p3803,p3804,p3805,p3806,p3807,p3808,p3809,p3810,p3811,p3812,p3813,p3814,p3815,p3816,p3817,p3818,p3819,p3820,p3821,p3822,p3823,p3824,p3825,p3826,p3827,p3828,p3829,p3830,p3831,p3832,p3833,p3834,p3835,p3836,p3837,p3838,p3839,p3840,p3841,p3842,p3843,p3844,p3845,p3846,p3847,p3848,p3849,p3850,p3851,p3852,p3853,p3854,p3855,p3856,p3857,p3858,p3859,p3860,p3861,p3862,p3863,p3864,p3865,p3866,p3867,p3868,p3869,p3870,p3871,p3872,p3873,p3874,p3875,p3876,p3877,p3878,p3879,p3880,p3881,p3882,p3883,p3884,p3885,p3886,p3887,p3888,p3889,p3890,p3891,p3892,p3893,p3894,p3895,p3896,p3897,p3898,p3899,p3900,p3901,p3902,p3903,p3904,p3905,p3906,p3907,p3908,p3909,p3910,p3911,p3912,p3913,p3914,p3915,p3916,p3917,p3918,p3919,p3920,p3921,p3922,p3923,p3924,p3925,p3926,p3927,p3928,p3929,p3930,p3931,p3932,p3933,p3934,p3935,p3936,p3937,p3938,p3939,p3940,p3941,p3942,p3943,p3944,p3945,p3946,p3947,p3948,p3949,p3950,p3951,p3952,p3953,p3954,p3955,p3956,p3957,p3958,p3959,p3960,p3961,p3962,p3963,p3964,p3965,p3966,p3967,p3968,p3969,p3970,p3971,p3972,p3973,p3974,p3975,p3976,p3977,p3978,p3979,p3980,p3981,p3982,p3983,p3984,p3985,p3986,p3987,p3988,p3989,p3990,p3991,p3992,p3993,p3994,p3995,p3996,p3997,p3998,p3999,p4000,p4001,p4002,p4003,p4004,p4005,p4006,p4007,p4008,p4009,p4010,p4011,p4012,p4013,p4014,p4015,p4016,p4017,p4018,p4019,p4020,p4021,p4022,p4023,p4024,p4025,p4026,p4027,p4028,p4029,p4030,p4031,p4032,p4033,p4034,p4035,p4036,p4037,p4038,p4039,p4040,p4041,p4042,p4043,p4044,p4045,p4046,p4047,p4048,p4049,p4050,p4051,p4052,p4053,p4054,p4055,p4056,p4057,p4058,p4059,p4060,p4061,p4062,p4063,p4064,p4065,p4066,p4067,p4068,p4069,p4070,p4071,p4072,p4073,p4074,p4075,p4076,p4077,p4078,p4079,p4080,p4081,p4082,p4083,p4084,p4085,p4086,p4087,p4088,p4089,p4090,p4091,p4092,p4093,p4094,p4095,p4096,p4097,p4098,p4099,p4100,p4101,p4102,p4103,p4104,p4105,p4106,p4107,p4108,p4109,p4110,p4111,p4112,p4113,p4114,p4115,p4116,p4117,p4118,p4119,p4120,p4121,p4122,p4123,p4124,p4125,p4126,p4127,p4128,p4129,p4130,p4131,p4132,p4133,p4134,p4135,p4136,p4137,p4138,p4139,p4140,p4141,p4142,p4143,p4144,p4145,p4146,p4147,p4148,p4149,p4150,p4151,p4152,p4153,p4154,p4155,p4156,p4157,p4158,p4159,p4160,p4161,p4162,p4163,p4164,p4165,p4166,p4167,p4168,p4169,p4170,p4171,p4172,p4173,p4174,p4175,p4176,p4177,p4178,p4179,p4180,p4181,p4182,p4183,p4184,p4185,p4186,p4187,p4188,p4189,p4190,p4191,p4192,p4193,p4194,p4195,p4196,p4197,p4198,p4199,p4200,p4201,p4202,p4203,p4204,p4205,p4206,p4207,p4208,p4209,p4210,p4211,p4212,p4213,p4214,p4215,p4216,p4217,p4218,p4219,p4220,p4221,p4222,p4223,p4224,p4225,p4226,p4227,p4228,p4229,p4230,p4231,p4232,p4233,p4234,p4235,p4236,p4237,p4238,p4239,p4240,p4241,p4242,p4243,p4244,p4245,p4246,p4247,p4248,p4249,p4250,p4251,p4252,p4253,p4254,p4255,p4256,p4257,p4258,p4259,p4260,p4261,p4262,p4263,p4264,p4265,p4266,p4267,p4268,p4269,p4270,p4271,p4272,p4273,p4274,p4275,p4276,p4277,p4278,p4279,p4280,p4281,p4282,p4283,p4284,p4285,p4286,p4287,p4288,p4289,p4290,p4291,p4292,p4293,p4294,p4295,p4296,p4297,p4298,p4299,p4300,p4301,p4302,p4303,p4304,p4305,p4306,p4307,p4308,p4309,p4310,p4311,p4312,p4313,p4314,p4315,p4316,p4317,p4318,p4319,p4320,p4321,p4322,p4323,p4324,p4325,p4326,p4327,p4328,p4329,p4330,p4331,p4332,p4333,p4334,p4335,p4336,p4337,p4338,p4339,p4340,p4341,p4342,p4343,p4344,p4345,p4346,p4347,p4348,p4349,p4350,p4351,p4352,p4353,p4354,p4355,p4356,p4357,p4358,p4359,p4360,p4361,p4362,p4363,p4364,p4365,p4366,p4367,p4368,p4369,p4370,p4371,p4372,p4373,p4374,p4375,p4376,p4377,p4378,p4379,p4380,p4381,p4382,p4383,p4384,p4385,p4386,p4387,p4388,p4389,p4390,p4391,p4392,p4393,p4394,p4395,p4396,p4397,p4398,p4399,p4400,p4401,p4402,p4403,p4404,p4405,p4406,p4407,p4408,p4409,p4410,p4411,p4412,p4413,p4414,p4415,p4416,p4417,p4418,p4419,p4420,p4421,p4422,p4423,p4424,p4425,p4426,p4427,p4428,p4429,p4430,p4431,p4432,p4433,p4434,p4435,p4436,p4437,p4438,p4439,p4440,p4441,p4442,p4443,p4444,p4445,p4446,p4447,p4448,p4449,p4450,p4451,p4452,p4453,p4454,p4455,p4456,p4457,p4458,p4459,p4460,p4461,p4462,p4463,p4464,p4465,p4466,p4467,p4468,p4469,p4470,p4471,p4472,p4473,p4474,p4475,p4476,p4477,p4478,p4479,p4480,p4481,p4482,p4483,p4484,p4485,p4486,p4487,p4488,p4489,p4490,p4491,p4492,p4493,p4494,p4495,p4496,p4497,p4498,p4499,p4500,p4501,p4502,p4503,p4504,p4505,p4506,p4507,p4508,p4509,p4510,p4511,p4512,p4513,p4514,p4515,p4516,p4517,p4518,p4519,p4520,p4521,p4522,p4523,p4524,p4525,p4526,p4527,p4528,p4529,p4530,p4531,p4532,p4533,p4534,p4535,p4536,p4537,p4538,p4539,p4540,p4541,p4542,p4543,p4544,p4545,p4546,p4547,p4548,p4549,p4550,p4551,p4552,p4553,p4554,p4555,p4556,p4557,p4558,p4559,p4560,p4561,p4562,p4563,p4564,p4565,p4566,p4567,p4568,p4569,p4570,p4571,p4572,p4573,p4574,p4575,p4576,p4577,p4578,p4579,p4580,p4581,p4582,p4583,p4584,p4585,p4586,p4587,p4588,p4589,p4590,p4591,p4592,p4593,p4594,p4595,p4596,p4597,p4598,p4599,p4600,p4601,p4602,p4603,p4604,p4605,p4606,p4607,p4608,p4609,p4610,p4611,p4612,p4613,p4614,p4615,p4616,p4617,p4618,p4619,p4620,p4621,p4622,p4623,p4624,p4625,p4626,p4627,p4628,p4629,p4630,p4631,p4632,p4633,p4634,p4635,p4636,p4637,p4638,p4639,p4640,p4641,p4642,p4643,p4644,p4645,p4646,p4647,p4648,p4649,p4650,p4651,p4652,p4653,p4654,p4655,p4656,p4657,p4658,p4659,p4660,p4661,p4662,p4663,p4664,p4665,p4666,p4667,p4668,p4669,p4670,p4671,p4672,p4673,p4674,p4675,p4676,p4677,p4678,p4679,p4680,p4681,p4682,p4683,p4684,p4685,p4686,p4687,p4688,p4689,p4690,p4691,p4692,p4693,p4694,p4695,p4696,p4697,p4698,p4699,p4700,p4701,p4702,p4703,p4704,p4705,p4706,p4707,p4708,p4709,p4710,p4711,p4712,p4713,p4714,p4715,p4716,p4717,p4718,p4719,p4720,p4721,p4722,p4723,p4724,p4725,p4726,p4727,p4728,p4729,p4730,p4731,p4732,p4733,p4734,p4735,p4736,p4737,p4738,p4739,p4740,p4741,p4742,p4743,p4744,p4745,p4746,p4747,p4748,p4749,p4750,p4751,p4752,p4753,p4754,p4755,p4756,p4757,p4758,p4759,p4760,p4761,p4762,p4763,p4764,p4765,p4766,p4767,p4768,p4769,p4770,p4771,p4772,p4773,p4774,p4775,p4776,p4777,p4778,p4779,p4780,p4781,p4782,p4783,p4784,p4785,p4786,p4787,p4788,p4789,p4790,p4791,p4792,p4793,p4794,p4795,p4796,p4797,p4798,p4799,p4800,p4801,p4802,p4803,p4804,p4805,p4806,p4807,p4808,p4809,p4810,p4811,p4812,p4813,p4814,p4815,p4816,p4817,p4818,p4819,p4820,p4821,p4822,p4823,p4824,p4825,p4826,p4827,p4828,p4829,p4830,p4831,p4832,p4833,p4834,p4835,p4836,p4837,p4838,p4839,p4840,p4841,p4842,p4843,p4844,p4845,p4846,p4847,p4848,p4849,p4850,p4851,p4852,p4853,p4854,p4855,p4856,p4857,p4858,p4859,p4860,p4861,p4862,p4863,p4864,p4865,p4866,p4867,p4868,p4869,p4870,p4871,p4872,p4873,p4874,p4875,p4876,p4877,p4878,p4879,p4880,p4881,p4882,p4883,p4884,p4885,p4886,p4887,p4888,p4889,p4890,p4891,p4892,p4893,p4894,p4895,p4896,p4897,p4898,p4899,p4900,p4901,p4902,p4903,p4904,p4905,p4906,p4907,p4908,p4909,p4910,p4911,p4912,p4913,p4914,p4915,p4916,p4917,p4918,p4919,p4920,p4921,p4922,p4923,p4924,p4925,p4926,p4927,p4928,p4929,p4930,p4931,p4932,p4933,p4934,p4935,p4936,p4937,p4938,p4939,p4940,p4941,p4942,p4943,p4944,p4945,p4946,p4947,p4948,p4949,p4950,p4951,p4952,p4953,p4954,p4955,p4956,p4957,p4958,p4959,p4960,p4961,p4962,p4963,p4964,p4965,p4966,p4967,p4968,p4969,p4970,p4971,p4972,p4973,p4974,p4975,p4976,p4977,p4978,p4979,p4980,p4981,p4982,p4983,p4984,p4985,p4986,p4987,p4988,p4989,p4990,p4991,p4992,p4993,p4994,p4995,p4996,p4997,p4998,p4999,p5000,p5001,p5002,p5003,p5004,p5005,p5006,p5007,p5008,p5009,p5010,p5011,p5012,p5013,p5014,p5015,p5016,p5017,p5018,p5019,p5020,p5021,p5022,p5023,p5024,p5025,p5026,p5027,p5028,p5029,p5030,p5031,p5032,p5033,p5034,p5035,p5036,p5037,p5038,p5039,p5040,p5041,p5042,p5043,p5044,p5045,p5046,p5047,p5048,p5049,p5050,p5051,p5052,p5053,p5054,p5055,p5056,p5057,p5058,p5059,p5060,p5061,p5062,p5063,p5064,p5065,p5066,p5067,p5068,p5069,p5070,p5071,p5072,p5073,p5074,p5075,p5076,p5077,p5078,p5079,p5080,p5081,p5082,p5083,p5084,p5085,p5086,p5087,p5088,p5089,p5090,p5091,p5092,p5093,p5094,p5095,p5096,p5097,p5098,p5099,p5100,p5101,p5102,p5103,p5104,p5105,p5106,p5107,p5108,p5109,p5110,p5111,p5112,p5113,p5114,p5115,p5116,p5117,p5118,p5119,p5120,p5121,p5122,p5123,p5124,p5125,p5126,p5127,p5128,p5129,p5130,p5131,p5132,p5133,p5134,p5135,p5136,p5137,p5138,p5139,p5140,p5141,p5142,p5143,p5144,p5145,p5146,p5147,p5148,p5149,p5150,p5151,p5152,p5153,p5154,p5155,p5156,p5157,p5158,p5159,p5160,p5161,p5162,p5163,p5164,p5165,p5166,p5167,p5168,p5169,p5170,p5171,p5172,p5173,p5174,p5175,p5176,p5177,p5178,p5179,p5180,p5181,p5182,p5183,p5184,p5185,p5186,p5187,p5188,p5189,p5190,p5191,p5192,p5193,p5194,p5195,p5196,p5197,p5198,p5199,p5200,p5201,p5202,p5203,p5204,p5205,p5206,p5207,p5208,p5209,p5210,p5211,p5212,p5213,p5214,p5215,p5216,p5217,p5218,p5219,p5220,p5221,p5222,p5223,p5224,p5225,p5226,p5227,p5228,p5229,p5230,p5231,p5232,p5233,p5234,p5235,p5236,p5237,p5238,p5239,p5240,p5241,p5242,p5243,p5244,p5245,p5246,p5247,p5248,p5249,p5250,p5251,p5252,p5253,p5254,p5255,p5256,p5257,p5258,p5259,p5260,p5261,p5262,p5263,p5264,p5265,p5266,p5267,p5268,p5269,p5270,p5271,p5272,p5273,p5274,p5275,p5276,p5277,p5278,p5279,p5280,p5281,p5282,p5283,p5284,p5285,p5286,p5287,p5288,p5289,p5290,p5291,p5292,p5293,p5294,p5295,p5296,p5297,p5298,p5299,p5300,p5301,p5302,p5303,p5304,p5305,p5306,p5307,p5308,p5309,p5310,p5311,p5312,p5313,p5314,p5315,p5316,p5317,p5318,p5319,p5320,p5321,p5322,p5323,p5324,p5325,p5326,p5327,p5328,p5329,p5330,p5331,p5332,p5333,p5334,p5335,p5336,p5337,p5338,p5339,p5340,p5341,p5342,p5343,p5344,p5345,p5346,p5347,p5348,p5349,p5350,p5351,p5352,p5353,p5354,p5355,p5356,p5357,p5358,p5359,p5360,p5361,p5362,p5363,p5364,p5365,p5366,p5367,p5368,p5369,p5370,p5371,p5372,p5373,p5374,p5375,p5376,p5377,p5378,p5379,p5380,p5381,p5382,p5383,p5384,p5385,p5386,p5387,p5388,p5389,p5390,p5391,p5392,p5393,p5394,p5395,p5396,p5397,p5398,p5399,p5400,p5401,p5402,p5403,p5404,p5405,p5406,p5407,p5408,p5409,p5410,p5411,p5412,p5413,p5414,p5415,p5416,p5417,p5418,p5419,p5420,p5421,p5422,p5423,p5424,p5425,p5426,p5427,p5428,p5429,p5430,p5431,p5432,p5433,p5434,p5435,p5436,p5437,p5438,p5439,p5440,p5441,p5442,p5443,p5444,p5445,p5446,p5447,p5448,p5449,p5450,p5451,p5452,p5453,p5454,p5455,p5456,p5457,p5458,p5459,p5460,p5461,p5462,p5463,p5464,p5465,p5466,p5467,p5468,p5469,p5470,p5471,p5472,p5473,p5474,p5475,p5476,p5477,p5478,p5479,p5480,p5481,p5482,p5483,p5484,p5485,p5486,p5487,p5488,p5489,p5490,p5491,p5492,p5493,p5494,p5495,p5496,p5497,p5498,p5499,p5500,p5501,p5502,p5503,p5504,p5505,p5506,p5507,p5508,p5509,p5510,p5511,p5512,p5513,p5514,p5515,p5516,p5517,p5518,p5519,p5520,p5521,p5522,p5523,p5524,p5525,p5526,p5527,p5528,p5529,p5530,p5531,p5532,p5533,p5534,p5535,p5536,p5537,p5538,p5539,p5540,p5541,p5542,p5543,p5544,p5545,p5546,p5547,p5548,p5549,p5550,p5551,p5552,p5553,p5554,p5555,p5556,p5557,p5558,p5559,p5560,p5561,p5562,p5563,p5564,p5565,p5566,p5567,p5568,p5569,p5570,p5571,p5572,p5573,p5574,p5575,p5576,p5577,p5578,p5579,p5580,p5581,p5582,p5583,p5584,p5585,p5586,p5587,p5588,p5589,p5590,p5591,p5592,p5593,p5594,p5595,p5596,p5597,p5598,p5599,p5600,p5601,p5602,p5603,p5604,p5605,p5606,p5607,p5608,p5609,p5610,p5611,p5612,p5613,p5614,p5615,p5616,p5617,p5618,p5619,p5620,p5621,p5622,p5623,p5624,p5625,p5626,p5627,p5628,p5629,p5630,p5631,p5632,p5633,p5634,p5635,p5636,p5637,p5638,p5639,p5640,p5641,p5642,p5643,p5644,p5645,p5646,p5647,p5648,p5649,p5650,p5651,p5652,p5653,p5654,p5655,p5656,p5657,p5658,p5659,p5660,p5661,p5662,p5663,p5664,p5665,p5666,p5667,p5668,p5669,p5670,p5671,p5672,p5673,p5674,p5675,p5676,p5677,p5678,p5679,p5680,p5681,p5682,p5683,p5684,p5685,p5686,p5687,p5688,p5689,p5690,p5691,p5692,p5693,p5694,p5695,p5696,p5697,p5698,p5699,p5700,p5701,p5702,p5703,p5704,p5705,p5706,p5707,p5708,p5709,p5710,p5711,p5712,p5713,p5714,p5715,p5716,p5717,p5718,p5719,p5720,p5721,p5722,p5723,p5724,p5725,p5726,p5727,p5728,p5729,p5730,p5731,p5732,p5733,p5734,p5735,p5736,p5737,p5738,p5739,p5740,p5741,p5742,p5743,p5744,p5745,p5746,p5747,p5748,p5749,p5750,p5751,p5752,p5753,p5754,p5755,p5756,p5757,p5758,p5759,p5760,p5761,p5762,p5763,p5764,p5765,p5766,p5767,p5768,p5769,p5770,p5771,p5772,p5773,p5774,p5775,p5776,p5777,p5778,p5779,p5780,p5781,p5782,p5783,p5784,p5785,p5786,p5787,p5788,p5789,p5790,p5791,p5792,p5793,p5794,p5795,p5796,p5797,p5798,p5799,p5800,p5801,p5802,p5803,p5804,p5805,p5806,p5807,p5808,p5809,p5810,p5811,p5812,p5813,p5814,p5815,p5816,p5817,p5818,p5819,p5820,p5821,p5822,p5823,p5824,p5825,p5826,p5827,p5828,p5829,p5830,p5831,p5832,p5833,p5834,p5835,p5836,p5837,p5838,p5839,p5840,p5841,p5842,p5843,p5844,p5845,p5846,p5847,p5848,p5849,p5850,p5851,p5852,p5853,p5854,p5855,p5856,p5857,p5858,p5859,p5860,p5861,p5862,p5863,p5864,p5865,p5866,p5867,p5868,p5869,p5870,p5871,p5872,p5873,p5874,p5875,p5876,p5877,p5878,p5879,p5880,p5881,p5882,p5883,p5884,p5885,p5886,p5887,p5888,p5889,p5890,p5891,p5892,p5893,p5894,p5895,p5896,p5897,p5898,p5899,p5900,p5901,p5902,p5903,p5904,p5905,p5906,p5907,p5908,p5909,p5910,p5911,p5912,p5913,p5914,p5915,p5916,p5917,p5918,p5919,p5920,p5921,p5922,p5923,p5924,p5925,p5926,p5927,p5928,p5929,p5930,p5931,p5932,p5933,p5934,p5935,p5936,p5937,p5938,p5939,p5940,p5941,p5942,p5943,p5944,p5945,p5946,p5947,p5948,p5949,p5950,p5951,p5952,p5953,p5954,p5955,p5956,p5957,p5958,p5959,p5960,p5961,p5962,p5963,p5964,p5965,p5966,p5967,p5968,p5969,p5970,p5971,p5972,p5973,p5974,p5975,p5976,p5977,p5978,p5979,p5980,p5981,p5982,p5983,p5984,p5985,p5986,p5987,p5988,p5989,p5990,p5991,p5992,p5993,p5994,p5995,p5996,p5997,p5998,p5999,p6000,p6001,p6002,p6003,p6004,p6005,p6006,p6007,p6008,p6009,p6010,p6011,p6012,p6013,p6014,p6015,p6016,p6017,p6018,p6019,p6020,p6021,p6022,p6023,p6024,p6025,p6026,p6027,p6028,p6029,p6030,p6031,p6032,p6033,p6034,p6035,p6036,p6037,p6038,p6039,p6040,p6041,p6042,p6043,p6044,p6045,p6046,p6047,p6048,p6049,p6050,p6051,p6052,p6053,p6054,p6055,p6056,p6057,p6058,p6059,p6060,p6061,p6062,p6063,p6064,p6065,p6066,p6067,p6068,p6069,p6070,p6071,p6072,p6073,p6074,p6075,p6076,p6077,p6078,p6079,p6080,p6081,p6082,p6083,p6084,p6085,p6086,p6087,p6088,p6089,p6090,p6091,p6092,p6093,p6094,p6095,p6096,p6097,p6098,p6099,p6100,p6101,p6102,p6103,p6104,p6105,p6106,p6107,p6108,p6109,p6110,p6111,p6112,p6113,p6114,p6115,p6116,p6117,p6118,p6119,p6120,p6121,p6122,p6123,p6124,p6125,p6126,p6127,p6128,p6129,p6130,p6131,p6132,p6133,p6134,p6135,p6136,p6137,p6138,p6139,p6140,p6141,p6142,p6143,p6144,p6145,p6146,p6147,p6148,p6149,p6150,p6151,p6152,p6153,p6154,p6155,p6156,p6157,p6158,p6159,p6160,p6161,p6162,p6163,p6164,p6165,p6166,p6167,p6168,p6169,p6170,p6171,p6172,p6173,p6174,p6175,p6176,p6177,p6178,p6179,p6180,p6181,p6182,p6183,p6184,p6185,p6186,p6187,p6188,p6189,p6190,p6191,p6192,p6193,p6194,p6195,p6196,p6197,p6198,p6199,p6200,p6201,p6202,p6203,p6204,p6205,p6206,p6207,p6208,p6209,p6210,p6211,p6212,p6213,p6214,p6215,p6216,p6217,p6218,p6219,p6220,p6221,p6222,p6223,p6224,p6225,p6226,p6227,p6228,p6229,p6230,p6231,p6232,p6233,p6234,p6235,p6236,p6237,p6238,p6239,p6240,p6241,p6242,p6243,p6244,p6245,p6246,p6247,p6248,p6249,p6250,p6251,p6252,p6253,p6254,p6255,p6256,p6257,p6258,p6259,p6260,p6261,p6262,p6263,p6264,p6265,p6266,p6267,p6268,p6269,p6270,p6271,p6272,p6273,p6274,p6275,p6276,p6277,p6278,p6279,p6280,p6281,p6282,p6283,p6284,p6285,p6286,p6287,p6288,p6289,p6290,p6291,p6292,p6293,p6294,p6295,p6296,p6297,p6298,p6299,p6300,p6301,p6302,p6303,p6304,p6305,p6306,p6307,p6308,p6309,p6310,p6311,p6312,p6313,p6314,p6315,p6316,p6317,p6318,p6319,p6320,p6321,p6322,p6323,p6324,p6325,p6326,p6327,p6328,p6329,p6330,p6331,p6332,p6333,p6334,p6335,p6336,p6337,p6338,p6339,p6340,p6341,p6342,p6343,p6344,p6345,p6346,p6347,p6348,p6349,p6350,p6351,p6352,p6353,p6354,p6355,p6356,p6357,p6358,p6359,p6360,p6361,p6362,p6363,p6364,p6365,p6366,p6367,p6368,p6369,p6370,p6371,p6372,p6373,p6374,p6375,p6376,p6377,p6378,p6379,p6380,p6381,p6382,p6383,p6384,p6385,p6386,p6387,p6388,p6389,p6390,p6391,p6392,p6393,p6394,p6395,p6396,p6397,p6398,p6399,p6400,p6401,p6402,p6403,p6404,p6405,p6406,p6407,p6408,p6409,p6410,p6411,p6412,p6413,p6414,p6415,p6416,p6417,p6418,p6419,p6420,p6421,p6422,p6423,p6424,p6425,p6426,p6427,p6428,p6429,p6430,p6431,p6432,p6433,p6434,p6435,p6436,p6437,p6438,p6439,p6440,p6441,p6442,p6443,p6444,p6445,p6446,p6447,p6448,p6449,p6450,p6451,p6452,p6453,p6454,p6455,p6456,p6457,p6458,p6459,p6460,p6461,p6462,p6463,p6464,p6465,p6466,p6467,p6468,p6469,p6470,p6471,p6472,p6473,p6474,p6475,p6476,p6477,p6478,p6479,p6480,p6481,p6482,p6483,p6484,p6485,p6486,p6487,p6488,p6489,p6490,p6491,p6492,p6493,p6494,p6495,p6496,p6497,p6498,p6499,p6500,p6501,p6502,p6503,p6504,p6505,p6506,p6507,p6508,p6509,p6510,p6511,p6512,p6513,p6514,p6515,p6516,p6517,p6518,p6519,p6520,p6521,p6522,p6523,p6524,p6525,p6526,p6527,p6528,p6529,p6530,p6531,p6532,p6533,p6534,p6535,p6536,p6537,p6538,p6539,p6540,p6541,p6542,p6543,p6544,p6545,p6546,p6547,p6548,p6549,p6550,p6551,p6552,p6553,p6554,p6555,p6556,p6557,p6558,p6559,p6560,p6561,p6562,p6563,p6564,p6565,p6566,p6567,p6568,p6569,p6570,p6571,p6572,p6573,p6574,p6575,p6576,p6577,p6578,p6579,p6580,p6581,p6582,p6583,p6584,p6585,p6586,p6587,p6588,p6589,p6590,p6591,p6592,p6593,p6594,p6595,p6596,p6597,p6598,p6599,p6600,p6601,p6602,p6603,p6604,p6605,p6606,p6607,p6608,p6609,p6610,p6611,p6612,p6613,p6614,p6615,p6616,p6617,p6618,p6619,p6620,p6621,p6622,p6623,p6624,p6625,p6626,p6627,p6628,p6629,p6630,p6631,p6632,p6633,p6634,p6635,p6636,p6637,p6638,p6639,p6640,p6641,p6642,p6643,p6644,p6645,p6646,p6647,p6648,p6649,p6650,p6651,p6652,p6653,p6654,p6655,p6656,p6657,p6658,p6659,p6660,p6661,p6662,p6663,p6664,p6665,p6666,p6667,p6668,p6669,p6670,p6671,p6672,p6673,p6674,p6675,p6676,p6677,p6678,p6679,p6680,p6681,p6682,p6683,p6684,p6685,p6686,p6687,p6688,p6689,p6690,p6691,p6692,p6693,p6694,p6695,p6696,p6697,p6698,p6699,p6700,p6701,p6702,p6703,p6704,p6705,p6706,p6707,p6708,p6709,p6710,p6711,p6712,p6713,p6714,p6715,p6716,p6717,p6718,p6719,p6720,p6721,p6722,p6723,p6724,p6725,p6726,p6727,p6728,p6729,p6730,p6731,p6732,p6733,p6734,p6735,p6736,p6737,p6738,p6739,p6740,p6741,p6742,p6743,p6744,p6745,p6746,p6747,p6748,p6749,p6750,p6751,p6752,p6753,p6754,p6755,p6756,p6757,p6758,p6759,p6760,p6761,p6762,p6763,p6764,p6765,p6766,p6767,p6768,p6769,p6770,p6771,p6772,p6773,p6774,p6775,p6776,p6777,p6778,p6779,p6780,p6781,p6782,p6783,p6784,p6785,p6786,p6787,p6788,p6789,p6790,p6791,p6792,p6793,p6794,p6795,p6796,p6797,p6798,p6799,p6800,p6801,p6802,p6803,p6804,p6805,p6806,p6807,p6808,p6809,p6810,p6811,p6812,p6813,p6814,p6815,p6816,p6817,p6818,p6819,p6820,p6821,p6822,p6823,p6824,p6825,p6826,p6827,p6828,p6829,p6830,p6831,p6832,p6833,p6834,p6835,p6836,p6837,p6838,p6839,p6840,p6841,p6842,p6843,p6844,p6845,p6846,p6847,p6848,p6849,p6850,p6851,p6852,p6853,p6854,p6855,p6856,p6857,p6858,p6859,p6860,p6861,p6862,p6863,p6864,p6865,p6866,p6867,p6868,p6869,p6870,p6871,p6872,p6873,p6874,p6875,p6876,p6877,p6878,p6879,p6880,p6881,p6882,p6883,p6884,p6885,p6886,p6887,p6888,p6889,p6890,p6891,p6892,p6893,p6894,p6895,p6896,p6897,p6898,p6899,p6900,p6901,p6902,p6903,p6904,p6905,p6906,p6907,p6908,p6909,p6910,p6911,p6912,p6913,p6914,p6915,p6916,p6917,p6918,p6919,p6920,p6921,p6922,p6923,p6924,p6925,p6926,p6927,p6928,p6929,p6930,p6931,p6932,p6933,p6934,p6935,p6936,p6937,p6938,p6939,p6940,p6941,p6942,p6943,p6944,p6945,p6946,p6947,p6948,p6949,p6950,p6951,p6952,p6953,p6954,p6955,p6956,p6957,p6958,p6959,p6960,p6961,p6962,p6963,p6964,p6965,p6966,p6967,p6968,p6969,p6970,p6971,p6972,p6973,p6974,p6975,p6976,p6977,p6978,p6979,p6980,p6981,p6982,p6983,p6984,p6985,p6986,p6987,p6988,p6989,p6990,p6991,p6992,p6993,p6994,p6995,p6996,p6997,p6998,p6999,p7000,p7001,p7002,p7003,p7004,p7005,p7006,p7007,p7008,p7009,p7010,p7011,p7012,p7013,p7014,p7015,p7016,p7017,p7018,p7019,p7020,p7021,p7022,p7023,p7024,p7025,p7026,p7027,p7028,p7029,p7030,p7031,p7032,p7033,p7034,p7035,p7036,p7037,p7038,p7039,p7040,p7041,p7042,p7043,p7044,p7045,p7046,p7047,p7048,p7049,p7050,p7051,p7052,p7053,p7054,p7055,p7056,p7057,p7058,p7059,p7060,p7061,p7062,p7063,p7064,p7065,p7066,p7067,p7068,p7069,p7070,p7071,p7072,p7073,p7074,p7075,p7076,p7077,p7078,p7079,p7080,p7081,p7082,p7083,p7084,p7085,p7086,p7087,p7088,p7089,p7090,p7091,p7092,p7093,p7094,p7095,p7096,p7097,p7098,p7099,p7100,p7101,p7102,p7103,p7104,p7105,p7106,p7107,p7108,p7109,p7110,p7111,p7112,p7113,p7114,p7115,p7116,p7117,p7118,p7119,p7120,p7121,p7122,p7123,p7124,p7125,p7126,p7127,p7128,p7129,p7130,p7131,p7132,p7133,p7134,p7135,p7136,p7137,p7138,p7139,p7140,p7141,p7142,p7143,p7144,p7145,p7146,p7147,p7148,p7149,p7150,p7151,p7152,p7153,p7154,p7155,p7156,p7157,p7158,p7159,p7160,p7161,p7162,p7163,p7164,p7165,p7166,p7167,p7168,p7169,p7170,p7171,p7172,p7173,p7174,p7175,p7176,p7177,p7178,p7179,p7180,p7181,p7182,p7183,p7184,p7185,p7186,p7187,p7188,p7189,p7190,p7191,p7192,p7193,p7194,p7195,p7196,p7197,p7198,p7199,p7200,p7201,p7202,p7203,p7204,p7205,p7206,p7207,p7208,p7209,p7210,p7211,p7212,p7213,p7214,p7215,p7216,p7217,p7218,p7219,p7220,p7221,p7222,p7223,p7224,p7225,p7226,p7227,p7228,p7229,p7230,p7231,p7232,p7233,p7234,p7235,p7236,p7237,p7238,p7239,p7240,p7241,p7242,p7243,p7244,p7245,p7246,p7247,p7248,p7249,p7250,p7251,p7252,p7253,p7254,p7255,p7256,p7257,p7258,p7259,p7260,p7261,p7262,p7263,p7264,p7265,p7266,p7267,p7268,p7269,p7270,p7271,p7272,p7273,p7274,p7275,p7276,p7277,p7278,p7279,p7280,p7281,p7282,p7283,p7284,p7285,p7286,p7287,p7288,p7289,p7290,p7291,p7292,p7293,p7294,p7295,p7296,p7297,p7298,p7299,p7300,p7301,p7302,p7303,p7304,p7305,p7306,p7307,p7308,p7309,p7310,p7311,p7312,p7313,p7314,p7315,p7316,p7317,p7318,p7319,p7320,p7321,p7322,p7323,p7324,p7325,p7326,p7327,p7328,p7329,p7330,p7331,p7332,p7333,p7334,p7335,p7336,p7337,p7338,p7339,p7340,p7341,p7342,p7343,p7344,p7345,p7346,p7347,p7348,p7349,p7350,p7351,p7352,p7353,p7354,p7355,p7356,p7357,p7358,p7359,p7360,p7361,p7362,p7363,p7364,p7365,p7366,p7367,p7368,p7369,p7370,p7371,p7372,p7373,p7374,p7375,p7376,p7377,p7378,p7379,p7380,p7381,p7382,p7383,p7384,p7385,p7386,p7387,p7388,p7389,p7390,p7391,p7392,p7393,p7394,p7395,p7396,p7397,p7398,p7399,p7400,p7401,p7402,p7403,p7404,p7405,p7406,p7407,p7408,p7409,p7410,p7411,p7412,p7413,p7414,p7415,p7416,p7417,p7418,p7419,p7420,p7421,p7422,p7423,p7424,p7425,p7426,p7427,p7428,p7429,p7430,p7431,p7432,p7433,p7434,p7435,p7436,p7437,p7438,p7439,p7440,p7441,p7442,p7443,p7444,p7445,p7446,p7447,p7448,p7449,p7450,p7451,p7452,p7453,p7454,p7455,p7456,p7457,p7458,p7459,p7460,p7461,p7462,p7463,p7464,p7465,p7466,p7467,p7468,p7469,p7470,p7471,p7472,p7473,p7474,p7475,p7476,p7477,p7478,p7479,p7480,p7481,p7482,p7483,p7484,p7485,p7486,p7487,p7488,p7489,p7490,p7491,p7492,p7493,p7494,p7495,p7496,p7497,p7498,p7499,p7500,p7501,p7502,p7503,p7504,p7505,p7506,p7507,p7508,p7509,p7510,p7511,p7512,p7513,p7514,p7515,p7516,p7517,p7518,p7519,p7520,p7521,p7522,p7523,p7524,p7525,p7526,p7527,p7528,p7529,p7530,p7531,p7532,p7533,p7534,p7535,p7536,p7537,p7538,p7539,p7540,p7541,p7542,p7543,p7544,p7545,p7546,p7547,p7548,p7549,p7550,p7551,p7552,p7553,p7554,p7555,p7556,p7557,p7558,p7559,p7560,p7561,p7562,p7563,p7564,p7565,p7566,p7567,p7568,p7569,p7570,p7571,p7572,p7573,p7574,p7575,p7576,p7577,p7578,p7579,p7580,p7581,p7582,p7583,p7584,p7585,p7586,p7587,p7588,p7589,p7590,p7591,p7592,p7593,p7594,p7595,p7596,p7597,p7598,p7599,p7600,p7601,p7602,p7603,p7604,p7605,p7606,p7607,p7608,p7609,p7610,p7611,p7612,p7613,p7614,p7615,p7616,p7617,p7618,p7619,p7620,p7621,p7622,p7623,p7624,p7625,p7626,p7627,p7628,p7629,p7630,p7631,p7632,p7633,p7634,p7635,p7636,p7637,p7638,p7639,p7640,p7641,p7642,p7643,p7644,p7645,p7646,p7647,p7648,p7649,p7650,p7651,p7652,p7653,p7654,p7655,p7656,p7657,p7658,p7659,p7660,p7661,p7662,p7663,p7664,p7665,p7666,p7667,p7668,p7669,p7670,p7671,p7672,p7673,p7674,p7675,p7676,p7677,p7678,p7679,p7680,p7681,p7682,p7683,p7684,p7685,p7686,p7687,p7688,p7689,p7690,p7691,p7692,p7693,p7694,p7695,p7696,p7697,p7698,p7699,p7700,p7701,p7702,p7703,p7704,p7705,p7706,p7707,p7708,p7709,p7710,p7711,p7712,p7713,p7714,p7715,p7716,p7717,p7718,p7719,p7720,p7721,p7722,p7723,p7724,p7725,p7726,p7727,p7728,p7729,p7730,p7731,p7732,p7733,p7734,p7735,p7736,p7737,p7738,p7739,p7740,p7741,p7742,p7743,p7744,p7745,p7746,p7747,p7748,p7749,p7750,p7751,p7752,p7753,p7754,p7755,p7756,p7757,p7758,p7759,p7760,p7761,p7762,p7763,p7764,p7765,p7766,p7767,p7768,p7769,p7770,p7771,p7772,p7773,p7774,p7775,p7776,p7777,p7778,p7779,p7780,p7781,p7782,p7783,p7784,p7785,p7786,p7787,p7788,p7789,p7790,p7791,p7792,p7793,p7794,p7795,p7796,p7797,p7798,p7799,p7800,p7801,p7802,p7803,p7804,p7805,p7806,p7807,p7808,p7809,p7810,p7811,p7812,p7813,p7814,p7815,p7816,p7817,p7818,p7819,p7820,p7821,p7822,p7823,p7824,p7825,p7826,p7827,p7828,p7829,p7830,p7831,p7832,p7833,p7834,p7835,p7836,p7837,p7838,p7839,p7840,p7841,p7842,p7843,p7844,p7845,p7846,p7847,p7848,p7849,p7850,p7851,p7852,p7853,p7854,p7855,p7856,p7857,p7858,p7859,p7860,p7861,p7862,p7863,p7864,p7865,p7866,p7867,p7868,p7869,p7870,p7871,p7872,p7873,p7874,p7875,p7876,p7877,p7878,p7879,p7880,p7881,p7882,p7883,p7884,p7885,p7886,p7887,p7888,p7889,p7890,p7891,p7892,p7893,p7894,p7895,p7896,p7897,p7898,p7899,p7900,p7901,p7902,p7903,p7904,p7905,p7906,p7907,p7908,p7909,p7910,p7911,p7912,p7913,p7914,p7915,p7916,p7917,p7918,p7919,p7920,p7921,p7922,p7923,p7924,p7925,p7926,p7927,p7928,p7929,p7930,p7931,p7932,p7933,p7934,p7935,p7936,p7937,p7938,p7939,p7940,p7941,p7942,p7943,p7944,p7945,p7946,p7947,p7948,p7949,p7950,p7951,p7952,p7953,p7954,p7955,p7956,p7957,p7958,p7959,p7960,p7961,p7962,p7963,p7964,p7965,p7966,p7967,p7968,p7969,p7970,p7971,p7972,p7973,p7974,p7975,p7976,p7977,p7978,p7979,p7980,p7981,p7982,p7983,p7984,p7985,p7986,p7987,p7988,p7989,p7990,p7991,p7992,p7993,p7994,p7995,p7996,p7997,p7998,p7999,p8000,p8001,p8002,p8003,p8004,p8005,p8006,p8007,p8008,p8009,p8010,p8011,p8012,p8013,p8014,p8015,p8016,p8017,p8018,p8019,p8020,p8021,p8022,p8023,p8024,p8025,p8026,p8027,p8028,p8029,p8030,p8031,p8032,p8033,p8034,p8035,p8036,p8037,p8038,p8039,p8040,p8041,p8042,p8043,p8044,p8045,p8046,p8047,p8048,p8049,p8050,p8051,p8052,p8053,p8054,p8055,p8056,p8057,p8058,p8059,p8060,p8061,p8062,p8063,p8064,p8065,p8066,p8067,p8068,p8069,p8070,p8071,p8072,p8073,p8074,p8075,p8076,p8077,p8078,p8079,p8080,p8081,p8082,p8083,p8084,p8085,p8086,p8087,p8088,p8089,p8090,p8091,p8092,p8093,p8094,p8095,p8096,p8097,p8098,p8099,p8100,p8101,p8102,p8103,p8104,p8105,p8106,p8107,p8108,p8109,p8110,p8111,p8112,p8113,p8114,p8115,p8116,p8117,p8118,p8119,p8120,p8121,p8122,p8123,p8124,p8125,p8126,p8127,p8128,p8129,p8130,p8131,p8132,p8133,p8134,p8135,p8136,p8137,p8138,p8139,p8140,p8141,p8142,p8143,p8144,p8145,p8146,p8147,p8148,p8149,p8150,p8151,p8152,p8153,p8154,p8155,p8156,p8157,p8158,p8159,p8160,p8161,p8162,p8163,p8164,p8165,p8166,p8167,p8168,p8169,p8170,p8171,p8172,p8173,p8174,p8175,p8176,p8177,p8178,p8179,p8180,p8181,p8182,p8183,p8184,p8185,p8186,p8187,p8188,p8189,p8190,p8191,p8192,p8193,p8194,p8195,p8196,p8197,p8198,p8199,p8200,p8201,p8202,p8203,p8204,p8205,p8206,p8207,p8208,p8209,p8210,p8211,p8212,p8213,p8214,p8215,p8216,p8217,p8218,p8219,p8220,p8221,p8222,p8223,p8224,p8225,p8226,p8227,p8228,p8229,p8230,p8231,p8232,p8233,p8234,p8235,p8236,p8237,p8238,p8239,p8240,p8241,p8242,p8243,p8244,p8245,p8246,p8247,p8248,p8249,p8250,p8251,p8252,p8253,p8254,p8255,p8256,p8257,p8258,p8259,p8260,p8261,p8262,p8263,p8264,p8265,p8266,p8267,p8268,p8269,p8270,p8271,p8272,p8273,p8274,p8275,p8276,p8277,p8278,p8279,p8280,p8281,p8282,p8283,p8284,p8285,p8286,p8287,p8288,p8289,p8290,p8291,p8292,p8293,p8294,p8295,p8296,p8297,p8298,p8299,p8300,p8301,p8302,p8303,p8304,p8305,p8306,p8307,p8308,p8309,p8310,p8311,p8312,p8313,p8314,p8315,p8316,p8317,p8318,p8319,p8320,p8321,p8322,p8323,p8324,p8325,p8326,p8327,p8328,p8329,p8330,p8331,p8332,p8333,p8334,p8335,p8336,p8337,p8338,p8339,p8340,p8341,p8342,p8343,p8344,p8345,p8346,p8347,p8348,p8349,p8350,p8351,p8352,p8353,p8354,p8355,p8356,p8357,p8358,p8359,p8360,p8361,p8362,p8363,p8364,p8365,p8366,p8367,p8368,p8369,p8370,p8371,p8372,p8373,p8374,p8375,p8376,p8377,p8378,p8379,p8380,p8381,p8382,p8383,p8384,p8385,p8386,p8387,p8388,p8389,p8390,p8391,p8392,p8393,p8394,p8395,p8396,p8397,p8398,p8399,p8400,p8401,p8402,p8403,p8404,p8405,p8406,p8407,p8408,p8409,p8410,p8411,p8412,p8413,p8414,p8415,p8416,p8417,p8418,p8419,p8420,p8421,p8422,p8423,p8424,p8425,p8426,p8427,p8428,p8429,p8430,p8431,p8432,p8433,p8434,p8435,p8436,p8437,p8438,p8439,p8440,p8441,p8442,p8443,p8444,p8445,p8446,p8447,p8448,p8449,p8450,p8451,p8452,p8453,p8454,p8455,p8456,p8457,p8458,p8459,p8460,p8461,p8462,p8463,p8464,p8465,p8466,p8467,p8468,p8469,p8470,p8471,p8472,p8473,p8474,p8475,p8476,p8477,p8478,p8479,p8480,p8481,p8482,p8483,p8484,p8485,p8486,p8487,p8488,p8489,p8490,p8491,p8492,p8493,p8494,p8495,p8496,p8497,p8498,p8499,p8500,p8501,p8502,p8503,p8504,p8505,p8506,p8507,p8508,p8509,p8510,p8511,p8512,p8513,p8514,p8515,p8516,p8517,p8518,p8519,p8520,p8521,p8522,p8523,p8524,p8525,p8526,p8527,p8528,p8529,p8530,p8531,p8532,p8533,p8534,p8535,p8536,p8537,p8538,p8539,p8540,p8541,p8542,p8543,p8544,p8545,p8546,p8547,p8548,p8549,p8550,p8551,p8552,p8553,p8554,p8555,p8556,p8557,p8558,p8559,p8560,p8561,p8562,p8563,p8564,p8565,p8566,p8567,p8568,p8569,p8570,p8571,p8572,p8573,p8574,p8575,p8576,p8577,p8578,p8579,p8580,p8581,p8582,p8583,p8584,p8585,p8586,p8587,p8588,p8589,p8590,p8591,p8592,p8593,p8594,p8595,p8596,p8597,p8598,p8599,p8600,p8601,p8602,p8603,p8604,p8605,p8606,p8607,p8608,p8609,p8610,p8611,p8612,p8613,p8614,p8615,p8616,p8617,p8618,p8619,p8620,p8621,p8622,p8623,p8624,p8625,p8626,p8627,p8628,p8629,p8630,p8631,p8632,p8633,p8634,p8635,p8636,p8637,p8638,p8639,p8640,p8641,p8642,p8643,p8644,p8645,p8646,p8647,p8648,p8649,p8650,p8651,p8652,p8653,p8654,p8655,p8656,p8657,p8658,p8659,p8660,p8661,p8662,p8663,p8664,p8665,p8666,p8667,p8668,p8669,p8670,p8671,p8672,p8673,p8674,p8675,p8676,p8677,p8678,p8679,p8680,p8681,p8682,p8683,p8684,p8685,p8686,p8687,p8688,p8689,p8690,p8691,p8692,p8693,p8694,p8695,p8696,p8697,p8698,p8699,p8700,p8701,p8702,p8703,p8704,p8705,p8706,p8707,p8708,p8709,p8710,p8711,p8712,p8713,p8714,p8715,p8716,p8717,p8718,p8719,p8720,p8721,p8722,p8723,p8724,p8725,p8726,p8727,p8728,p8729,p8730,p8731,p8732,p8733,p8734,p8735,p8736,p8737,p8738,p8739,p8740,p8741,p8742,p8743,p8744,p8745,p8746,p8747,p8748,p8749,p8750,p8751,p8752,p8753,p8754,p8755,p8756,p8757,p8758,p8759,p8760,p8761,p8762,p8763,p8764,p8765,p8766,p8767,p8768,p8769,p8770,p8771,p8772,p8773,p8774,p8775,p8776,p8777,p8778,p8779,p8780,p8781,p8782,p8783,p8784,p8785,p8786,p8787,p8788,p8789,p8790,p8791,p8792,p8793,p8794,p8795,p8796,p8797,p8798,p8799,p8800,p8801,p8802,p8803,p8804,p8805,p8806,p8807,p8808,p8809,p8810,p8811,p8812,p8813,p8814,p8815,p8816,p8817,p8818,p8819,p8820,p8821,p8822,p8823,p8824,p8825,p8826,p8827,p8828,p8829,p8830,p8831,p8832,p8833,p8834,p8835,p8836,p8837,p8838,p8839,p8840,p8841,p8842,p8843,p8844,p8845,p8846,p8847,p8848,p8849,p8850,p8851,p8852,p8853,p8854,p8855,p8856,p8857,p8858,p8859,p8860,p8861,p8862,p8863,p8864,p8865,p8866,p8867,p8868,p8869,p8870,p8871,p8872,p8873,p8874,p8875,p8876,p8877,p8878,p8879,p8880,p8881,p8882,p8883,p8884,p8885,p8886,p8887,p8888,p8889,p8890,p8891,p8892,p8893,p8894,p8895,p8896,p8897,p8898,p8899,p8900,p8901,p8902,p8903,p8904,p8905,p8906,p8907,p8908,p8909,p8910,p8911,p8912,p8913,p8914,p8915,p8916,p8917,p8918,p8919,p8920,p8921,p8922,p8923,p8924,p8925,p8926,p8927,p8928,p8929,p8930,p8931,p8932,p8933,p8934,p8935,p8936,p8937,p8938,p8939,p8940,p8941,p8942,p8943,p8944,p8945,p8946,p8947,p8948,p8949,p8950,p8951,p8952,p8953,p8954,p8955,p8956,p8957,p8958,p8959,p8960,p8961,p8962,p8963,p8964,p8965,p8966,p8967,p8968,p8969,p8970,p8971,p8972,p8973,p8974,p8975,p8976,p8977,p8978,p8979,p8980,p8981,p8982,p8983,p8984,p8985,p8986,p8987,p8988,p8989,p8990,p8991,p8992,p8993,p8994,p8995,p8996,p8997,p8998,p8999,p9000,p9001,p9002,p9003,p9004,p9005,p9006,p9007,p9008,p9009,p9010,p9011,p9012,p9013,p9014,p9015,p9016,p9017,p9018,p9019,p9020,p9021,p9022,p9023,p9024,p9025,p9026,p9027,p9028,p9029,p9030,p9031,p9032,p9033,p9034,p9035,p9036,p9037,p9038,p9039,p9040,p9041,p9042,p9043,p9044,p9045,p9046,p9047,p9048,p9049,p9050,p9051,p9052,p9053,p9054,p9055,p9056,p9057,p9058,p9059,p9060,p9061,p9062,p9063,p9064,p9065,p9066,p9067,p9068,p9069,p9070,p9071,p9072,p9073,p9074,p9075,p9076,p9077,p9078,p9079,p9080,p9081,p9082,p9083,p9084,p9085,p9086,p9087,p9088,p9089,p9090,p9091,p9092,p9093,p9094,p9095,p9096,p9097,p9098,p9099,p9100,p9101,p9102,p9103,p9104,p9105,p9106,p9107,p9108,p9109,p9110,p9111,p9112,p9113,p9114,p9115,p9116,p9117,p9118,p9119,p9120,p9121,p9122,p9123,p9124,p9125,p9126,p9127,p9128,p9129,p9130,p9131,p9132,p9133,p9134,p9135,p9136,p9137,p9138,p9139,p9140,p9141,p9142,p9143,p9144,p9145,p9146,p9147,p9148,p9149,p9150,p9151,p9152,p9153,p9154,p9155,p9156,p9157,p9158,p9159,p9160,p9161,p9162,p9163,p9164,p9165,p9166,p9167,p9168,p9169,p9170,p9171,p9172,p9173,p9174,p9175,p9176,p9177,p9178,p9179,p9180,p9181,p9182,p9183,p9184,p9185,p9186,p9187,p9188,p9189,p9190,p9191,p9192,p9193,p9194,p9195,p9196,p9197,p9198,p9199,p9200,p9201,p9202,p9203,p9204,p9205,p9206,p9207,p9208,p9209,p9210,p9211,p9212,p9213,p9214,p9215,p9216,p9217,p9218,p9219,p9220,p9221,p9222,p9223,p9224,p9225,p9226,p9227,p9228,p9229,p9230,p9231,p9232,p9233,p9234,p9235,p9236,p9237,p9238,p9239,p9240,p9241,p9242,p9243,p9244,p9245,p9246,p9247,p9248,p9249,p9250,p9251,p9252,p9253,p9254,p9255,p9256,p9257,p9258,p9259,p9260,p9261,p9262,p9263,p9264,p9265,p9266,p9267,p9268,p9269,p9270,p9271,p9272,p9273,p9274,p9275,p9276,p9277,p9278,p9279,p9280,p9281,p9282,p9283,p9284,p9285,p9286,p9287,p9288,p9289,p9290,p9291,p9292,p9293,p9294,p9295,p9296,p9297,p9298,p9299,p9300,p9301,p9302,p9303,p9304,p9305,p9306,p9307,p9308,p9309,p9310,p9311,p9312,p9313,p9314,p9315,p9316,p9317,p9318,p9319,p9320,p9321,p9322,p9323,p9324,p9325,p9326,p9327,p9328,p9329,p9330,p9331,p9332,p9333,p9334,p9335,p9336,p9337,p9338,p9339,p9340,p9341,p9342,p9343,p9344,p9345,p9346,p9347,p9348,p9349,p9350,p9351,p9352,p9353,p9354,p9355,p9356,p9357,p9358,p9359,p9360,p9361,p9362,p9363,p9364,p9365,p9366,p9367,p9368,p9369,p9370,p9371,p9372,p9373,p9374,p9375,p9376,p9377,p9378,p9379,p9380,p9381,p9382,p9383,p9384,p9385,p9386,p9387,p9388,p9389,p9390,p9391,p9392,p9393,p9394,p9395,p9396,p9397,p9398,p9399,p9400,p9401,p9402,p9403,p9404,p9405,p9406,p9407,p9408,p9409,p9410,p9411,p9412,p9413,p9414,p9415,p9416,p9417,p9418,p9419,p9420,p9421,p9422,p9423,p9424,p9425,p9426,p9427,p9428,p9429,p9430,p9431,p9432,p9433,p9434,p9435,p9436,p9437,p9438,p9439,p9440,p9441,p9442,p9443,p9444,p9445,p9446,p9447,p9448,p9449,p9450,p9451,p9452,p9453,p9454,p9455,p9456,p9457,p9458,p9459,p9460,p9461,p9462,p9463,p9464,p9465,p9466,p9467,p9468,p9469,p9470,p9471,p9472,p9473,p9474,p9475,p9476,p9477,p9478,p9479,p9480,p9481,p9482,p9483,p9484,p9485,p9486,p9487,p9488,p9489,p9490,p9491,p9492,p9493,p9494,p9495,p9496,p9497,p9498,p9499,p9500,p9501,p9502,p9503,p9504,p9505,p9506,p9507,p9508,p9509,p9510,p9511,p9512,p9513,p9514,p9515,p9516,p9517,p9518,p9519,p9520,p9521,p9522,p9523,p9524,p9525,p9526,p9527,p9528,p9529,p9530,p9531,p9532,p9533,p9534,p9535,p9536,p9537,p9538,p9539,p9540,p9541,p9542,p9543,p9544,p9545,p9546,p9547,p9548,p9549,p9550,p9551,p9552,p9553,p9554,p9555,p9556,p9557,p9558,p9559,p9560,p9561,p9562,p9563,p9564,p9565,p9566,p9567,p9568,p9569,p9570,p9571,p9572,p9573,p9574,p9575,p9576,p9577,p9578,p9579,p9580,p9581,p9582,p9583,p9584,p9585,p9586,p9587,p9588,p9589,p9590,p9591,p9592,p9593,p9594,p9595,p9596,p9597,p9598,p9599,p9600,p9601,p9602,p9603,p9604,p9605,p9606,p9607,p9608,p9609,p9610,p9611,p9612,p9613,p9614,p9615,p9616,p9617,p9618,p9619,p9620,p9621,p9622,p9623,p9624,p9625,p9626,p9627,p9628,p9629,p9630,p9631,p9632,p9633,p9634,p9635,p9636,p9637,p9638,p9639,p9640,p9641,p9642,p9643,p9644,p9645,p9646,p9647,p9648,p9649,p9650,p9651,p9652,p9653,p9654,p9655,p9656,p9657,p9658,p9659,p9660,p9661,p9662,p9663,p9664,p9665,p9666,p9667,p9668,p9669,p9670,p9671,p9672,p9673,p9674,p9675,p9676,p9677,p9678,p9679,p9680,p9681,p9682,p9683,p9684,p9685,p9686,p9687,p9688,p9689,p9690,p9691,p9692,p9693,p9694,p9695,p9696,p9697,p9698,p9699,p9700,p9701,p9702,p9703,p9704,p9705,p9706,p9707,p9708,p9709,p9710,p9711,p9712,p9713,p9714,p9715,p9716,p9717,p9718,p9719,p9720,p9721,p9722,p9723,p9724,p9725,p9726,p9727,p9728,p9729,p9730,p9731,p9732,p9733,p9734,p9735,p9736,p9737,p9738,p9739,p9740,p9741,p9742,p9743,p9744,p9745,p9746,p9747,p9748,p9749,p9750,p9751,p9752,p9753,p9754,p9755,p9756,p9757,p9758,p9759,p9760,p9761,p9762,p9763,p9764,p9765,p9766,p9767,p9768,p9769,p9770,p9771,p9772,p9773,p9774,p9775,p9776,p9777,p9778,p9779,p9780,p9781,p9782,p9783,p9784,p9785,p9786,p9787,p9788,p9789,p9790,p9791,p9792,p9793,p9794,p9795,p9796,p9797,p9798,p9799,p9800,p9801,p9802,p9803,p9804,p9805,p9806,p9807,p9808,p9809,p9810,p9811,p9812,p9813,p9814,p9815,p9816,p9817,p9818,p9819,p9820,p9821,p9822,p9823,p9824,p9825,p9826,p9827,p9828,p9829,p9830,p9831,p9832,p9833,p9834,p9835,p9836,p9837,p9838,p9839,p9840,p9841,p9842,p9843,p9844,p9845,p9846,p9847,p9848,p9849,p9850,p9851,p9852,p9853,p9854,p9855,p9856,p9857,p9858,p9859,p9860,p9861,p9862,p9863,p9864,p9865,p9866,p9867,p9868,p9869,p9870,p9871,p9872,p9873,p9874,p9875,p9876,p9877,p9878,p9879,p9880,p9881,p9882,p9883,p9884,p9885,p9886,p9887,p9888,p9889,p9890,p9891,p9892,p9893,p9894,p9895,p9896,p9897,p9898,p9899,p9900,p9901,p9902,p9903,p9904,p9905,p9906,p9907,p9908,p9909,p9910,p9911,p9912,p9913,p9914,p9915,p9916,p9917,p9918,p9919,p9920,p9921,p9922,p9923,p9924,p9925,p9926,p9927,p9928,p9929,p9930,p9931,p9932,p9933,p9934,p9935,p9936,p9937,p9938,p9939,p9940,p9941,p9942,p9943,p9944,p9945,p9946,p9947,p9948,p9949,p9950,p9951,p9952,p9953,p9954,p9955,p9956,p9957,p9958,p9959,p9960,p9961,p9962,p9963,p9964,p9965,p9966,p9967,p9968,p9969,p9970,p9971,p9972,p9973,p9974,p9975,p9976,p9977,p9978,p9979,p9980,p9981,p9982,p9983,p9984,p9985,p9986,p9987,p9988,p9989,p9990,p9991,p9992,p9993,p9994,p9995,p9996,p9997,p9998,p9999,p10000,p10001,p10002,p10003,p10004,p10005,p10006,p10007,p10008,p10009,p10010,p10011,p10012,p10013,p10014,p10015,p10016,p10017,p10018,p10019,p10020,p10021,p10022,p10023,p10024,p10025,p10026,p10027,p10028,p10029,p10030,p10031,p10032,p10033,p10034,p10035,p10036,p10037,p10038,p10039,p10040,p10041,p10042,p10043,p10044,p10045,p10046,p10047,p10048,p10049,p10050,p10051,p10052,p10053,p10054,p10055,p10056,p10057,p10058,p10059,p10060,p10061,p10062,p10063,p10064,p10065,p10066,p10067,p10068,p10069,p10070,p10071,p10072,p10073,p10074,p10075,p10076,p10077,p10078,p10079,p10080,p10081,p10082,p10083,p10084,p10085,p10086,p10087,p10088,p10089,p10090,p10091,p10092,p10093,p10094,p10095,p10096,p10097,p10098,p10099,p10100,p10101,p10102,p10103,p10104,p10105,p10106,p10107,p10108,p10109,p10110,p10111,p10112,p10113,p10114,p10115,p10116,p10117,p10118,p10119,p10120,p10121,p10122,p10123,p10124,p10125,p10126,p10127,p10128,p10129,p10130,p10131,p10132,p10133,p10134,p10135,p10136,p10137,p10138,p10139,p10140,p10141,p10142,p10143,p10144,p10145,p10146,p10147,p10148,p10149,p10150,p10151,p10152,p10153,p10154,p10155,p10156,p10157,p10158,p10159,p10160,p10161,p10162,p10163,p10164,p10165,p10166,p10167,p10168,p10169,p10170,p10171,p10172,p10173,p10174,p10175,p10176,p10177,p10178,p10179,p10180,p10181,p10182,p10183,p10184,p10185,p10186,p10187,p10188,p10189,p10190,p10191,p10192,p10193,p10194,p10195,p10196,p10197,p10198,p10199,p10200,p10201,p10202,p10203,p10204,p10205,p10206,p10207,p10208,p10209,p10210,p10211,p10212,p10213,p10214,p10215,p10216,p10217,p10218,p10219,p10220,p10221,p10222,p10223,p10224,p10225,p10226,p10227,p10228,p10229,p10230,p10231,p10232,p10233,p10234,p10235,p10236,p10237,p10238,p10239,p10240,p10241,p10242,p10243,p10244,p10245,p10246,p10247,p10248,p10249,p10250,p10251,p10252,p10253,p10254,p10255,p10256,p10257,p10258,p10259,p10260,p10261,p10262,p10263,p10264,p10265,p10266,p10267,p10268,p10269,p10270,p10271,p10272,p10273,p10274,p10275,p10276,p10277,p10278,p10279,p10280,p10281,p10282,p10283,p10284,p10285,p10286,p10287,p10288,p10289,p10290,p10291,p10292,p10293,p10294,p10295,p10296,p10297,p10298,p10299,p10300,p10301,p10302,p10303,p10304,p10305,p10306,p10307,p10308,p10309,p10310,p10311,p10312,p10313,p10314,p10315,p10316,p10317,p10318,p10319,p10320,p10321,p10322,p10323,p10324,p10325,p10326,p10327,p10328,p10329,p10330,p10331,p10332,p10333,p10334,p10335,p10336,p10337,p10338,p10339,p10340,p10341,p10342,p10343,p10344,p10345,p10346,p10347,p10348,p10349,p10350,p10351,p10352,p10353,p10354,p10355,p10356,p10357,p10358,p10359,p10360,p10361,p10362,p10363,p10364,p10365,p10366,p10367,p10368,p10369,p10370,p10371,p10372,p10373,p10374,p10375,p10376,p10377,p10378,p10379,p10380,p10381,p10382,p10383,p10384,p10385,p10386,p10387,p10388,p10389,p10390,p10391,p10392,p10393,p10394,p10395,p10396,p10397,p10398,p10399,p10400,p10401,p10402,p10403,p10404,p10405,p10406,p10407,p10408,p10409,p10410,p10411,p10412,p10413,p10414,p10415,p10416,p10417,p10418,p10419,p10420,p10421,p10422,p10423,p10424,p10425,p10426,p10427,p10428,p10429,p10430,p10431,p10432,p10433,p10434,p10435,p10436,p10437,p10438,p10439,p10440,p10441,p10442,p10443,p10444,p10445,p10446,p10447,p10448,p10449,p10450,p10451,p10452,p10453,p10454,p10455,p10456,p10457,p10458,p10459,p10460,p10461,p10462,p10463,p10464,p10465,p10466,p10467,p10468,p10469,p10470,p10471,p10472,p10473,p10474,p10475,p10476,p10477,p10478,p10479,p10480,p10481,p10482,p10483,p10484,p10485,p10486,p10487,p10488,p10489,p10490,p10491,p10492,p10493,p10494,p10495,p10496,p10497,p10498,p10499,p10500,p10501,p10502,p10503,p10504,p10505,p10506,p10507,p10508,p10509,p10510,p10511,p10512,p10513,p10514,p10515,p10516,p10517,p10518,p10519,p10520,p10521,p10522,p10523,p10524,p10525,p10526,p10527,p10528,p10529,p10530,p10531,p10532,p10533,p10534,p10535,p10536,p10537,p10538,p10539,p10540,p10541,p10542,p10543,p10544,p10545,p10546,p10547,p10548,p10549,p10550,p10551,p10552,p10553,p10554,p10555,p10556,p10557,p10558,p10559,p10560,p10561,p10562,p10563,p10564,p10565,p10566,p10567,p10568,p10569,p10570,p10571,p10572,p10573,p10574,p10575,p10576,p10577,p10578,p10579,p10580,p10581,p10582,p10583,p10584,p10585,p10586,p10587,p10588,p10589,p10590,p10591,p10592,p10593,p10594,p10595,p10596,p10597,p10598,p10599,p10600,p10601,p10602,p10603,p10604,p10605,p10606,p10607,p10608,p10609,p10610,p10611,p10612,p10613,p10614,p10615,p10616,p10617,p10618,p10619,p10620,p10621,p10622,p10623,p10624,p10625,p10626,p10627,p10628,p10629,p10630,p10631,p10632,p10633,p10634,p10635,p10636,p10637,p10638,p10639,p10640,p10641,p10642,p10643,p10644,p10645,p10646,p10647,p10648,p10649,p10650,p10651,p10652,p10653,p10654,p10655,p10656,p10657,p10658,p10659,p10660,p10661,p10662,p10663,p10664,p10665,p10666,p10667,p10668,p10669,p10670,p10671,p10672,p10673,p10674,p10675,p10676,p10677,p10678,p10679,p10680,p10681,p10682,p10683,p10684,p10685,p10686,p10687,p10688,p10689,p10690,p10691,p10692,p10693,p10694,p10695,p10696,p10697,p10698,p10699,p10700,p10701,p10702,p10703,p10704,p10705,p10706,p10707,p10708,p10709,p10710,p10711,p10712,p10713,p10714,p10715,p10716,p10717,p10718,p10719,p10720,p10721,p10722,p10723,p10724,p10725,p10726,p10727,p10728,p10729,p10730,p10731,p10732,p10733,p10734,p10735,p10736,p10737,p10738,p10739,p10740,p10741,p10742,p10743,p10744,p10745,p10746,p10747,p10748,p10749,p10750,p10751,p10752,p10753,p10754,p10755,p10756,p10757,p10758,p10759,p10760,p10761,p10762,p10763,p10764,p10765,p10766,p10767,p10768,p10769,p10770,p10771,p10772,p10773,p10774,p10775,p10776,p10777,p10778,p10779,p10780,p10781,p10782,p10783,p10784,p10785,p10786,p10787,p10788,p10789,p10790,p10791,p10792,p10793,p10794,p10795,p10796,p10797,p10798,p10799,p10800,p10801,p10802,p10803,p10804,p10805,p10806,p10807,p10808,p10809,p10810,p10811,p10812,p10813,p10814,p10815,p10816,p10817,p10818,p10819,p10820,p10821,p10822,p10823,p10824,p10825,p10826,p10827,p10828,p10829,p10830,p10831,p10832,p10833,p10834,p10835,p10836,p10837,p10838,p10839,p10840,p10841,p10842,p10843,p10844,p10845,p10846,p10847,p10848,p10849,p10850,p10851,p10852,p10853,p10854,p10855,p10856,p10857,p10858,p10859,p10860,p10861,p10862,p10863,p10864,p10865,p10866,p10867,p10868,p10869,p10870,p10871,p10872,p10873,p10874,p10875,p10876,p10877,p10878,p10879,p10880,p10881,p10882,p10883,p10884,p10885,p10886,p10887,p10888,p10889,p10890,p10891,p10892,p10893,p10894,p10895,p10896,p10897,p10898,p10899,p10900,p10901,p10902,p10903,p10904,p10905,p10906,p10907,p10908,p10909,p10910,p10911,p10912,p10913,p10914,p10915,p10916,p10917,p10918,p10919,p10920,p10921,p10922,p10923,p10924,p10925,p10926,p10927,p10928,p10929,p10930,p10931,p10932,p10933,p10934,p10935,p10936,p10937,p10938,p10939,p10940,p10941,p10942,p10943,p10944,p10945,p10946,p10947,p10948,p10949,p10950,p10951,p10952,p10953,p10954,p10955,p10956,p10957,p10958,p10959,p10960,p10961,p10962,p10963,p10964,p10965,p10966,p10967,p10968,p10969,p10970,p10971,p10972,p10973,p10974,p10975,p10976,p10977,p10978,p10979,p10980,p10981,p10982,p10983,p10984,p10985,p10986,p10987,p10988,p10989,p10990,p10991,p10992,p10993,p10994,p10995,p10996,p10997,p10998,p10999,p11000,p11001,p11002,p11003,p11004,p11005,p11006,p11007,p11008,p11009,p11010,p11011,p11012,p11013,p11014,p11015,p11016,p11017,p11018,p11019,p11020,p11021,p11022,p11023,p11024,p11025,p11026,p11027,p11028,p11029,p11030,p11031,p11032,p11033,p11034,p11035,p11036,p11037,p11038,p11039,p11040,p11041,p11042,p11043,p11044,p11045,p11046,p11047,p11048,p11049,p11050,p11051,p11052,p11053,p11054,p11055,p11056,p11057,p11058,p11059,p11060,p11061,p11062,p11063,p11064,p11065,p11066,p11067,p11068,p11069,p11070,p11071,p11072,p11073,p11074,p11075,p11076,p11077,p11078,p11079,p11080,p11081,p11082,p11083,p11084,p11085,p11086,p11087,p11088,p11089,p11090,p11091,p11092,p11093,p11094,p11095,p11096,p11097,p11098,p11099,p11100,p11101,p11102,p11103,p11104,p11105,p11106,p11107,p11108,p11109,p11110,p11111,p11112,p11113,p11114,p11115,p11116,p11117,p11118,p11119,p11120,p11121,p11122,p11123,p11124,p11125,p11126,p11127,p11128,p11129,p11130,p11131,p11132,p11133,p11134,p11135,p11136,p11137,p11138,p11139,p11140,p11141,p11142,p11143,p11144,p11145,p11146,p11147,p11148,p11149,p11150,p11151,p11152,p11153,p11154,p11155,p11156,p11157,p11158,p11159,p11160,p11161,p11162,p11163,p11164,p11165,p11166,p11167,p11168,p11169,p11170,p11171,p11172,p11173,p11174,p11175,p11176,p11177,p11178,p11179,p11180,p11181,p11182,p11183,p11184,p11185,p11186,p11187,p11188,p11189,p11190,p11191,p11192,p11193,p11194,p11195,p11196,p11197,p11198,p11199,p11200,p11201,p11202,p11203,p11204,p11205,p11206,p11207,p11208,p11209,p11210,p11211,p11212,p11213,p11214,p11215,p11216,p11217,p11218,p11219,p11220,p11221,p11222,p11223,p11224,p11225,p11226,p11227,p11228,p11229,p11230,p11231,p11232,p11233,p11234,p11235,p11236,p11237,p11238,p11239,p11240,p11241,p11242,p11243,p11244,p11245,p11246,p11247,p11248,p11249,p11250,p11251,p11252,p11253,p11254,p11255,p11256,p11257,p11258,p11259,p11260,p11261,p11262,p11263,p11264,p11265,p11266,p11267,p11268,p11269,p11270,p11271,p11272,p11273,p11274,p11275,p11276,p11277,p11278,p11279,p11280,p11281,p11282,p11283,p11284,p11285,p11286,p11287,p11288,p11289,p11290,p11291,p11292,p11293,p11294,p11295,p11296,p11297,p11298,p11299,p11300,p11301,p11302,p11303,p11304,p11305,p11306,p11307,p11308,p11309,p11310,p11311,p11312,p11313,p11314,p11315,p11316,p11317,p11318,p11319,p11320,p11321,p11322,p11323,p11324,p11325,p11326,p11327,p11328,p11329,p11330,p11331,p11332,p11333,p11334,p11335,p11336,p11337,p11338,p11339,p11340,p11341,p11342,p11343,p11344,p11345,p11346,p11347,p11348,p11349,p11350,p11351,p11352,p11353,p11354,p11355,p11356,p11357,p11358,p11359,p11360,p11361,p11362,p11363,p11364,p11365,p11366,p11367,p11368,p11369,p11370,p11371,p11372,p11373,p11374,p11375,p11376,p11377,p11378,p11379,p11380,p11381,p11382,p11383,p11384,p11385,p11386,p11387,p11388,p11389,p11390,p11391,p11392,p11393,p11394,p11395,p11396,p11397,p11398,p11399,p11400,p11401,p11402,p11403,p11404,p11405,p11406,p11407,p11408,p11409,p11410,p11411,p11412,p11413,p11414,p11415,p11416,p11417,p11418,p11419,p11420,p11421,p11422,p11423,p11424,p11425,p11426,p11427,p11428,p11429,p11430,p11431,p11432,p11433,p11434,p11435,p11436,p11437,p11438,p11439,p11440,p11441,p11442,p11443,p11444,p11445,p11446,p11447,p11448,p11449,p11450,p11451,p11452,p11453,p11454,p11455,p11456,p11457,p11458,p11459,p11460,p11461,p11462,p11463,p11464,p11465,p11466,p11467,p11468,p11469,p11470,p11471,p11472,p11473,p11474,p11475,p11476,p11477,p11478,p11479,p11480,p11481,p11482,p11483,p11484,p11485,p11486,p11487,p11488,p11489,p11490,p11491,p11492,p11493,p11494,p11495,p11496,p11497,p11498,p11499,p11500,p11501,p11502,p11503,p11504,p11505,p11506,p11507,p11508,p11509,p11510,p11511,p11512,p11513,p11514,p11515,p11516,p11517,p11518,p11519,p11520,p11521,p11522,p11523,p11524,p11525,p11526,p11527,p11528,p11529,p11530,p11531,p11532,p11533,p11534,p11535,p11536,p11537,p11538,p11539,p11540,p11541,p11542,p11543,p11544,p11545,p11546,p11547,p11548,p11549,p11550,p11551,p11552,p11553,p11554,p11555,p11556,p11557,p11558,p11559,p11560,p11561,p11562,p11563,p11564,p11565,p11566,p11567,p11568,p11569,p11570,p11571,p11572,p11573,p11574,p11575,p11576,p11577,p11578,p11579,p11580,p11581,p11582,p11583,p11584,p11585,p11586,p11587,p11588,p11589,p11590,p11591,p11592,p11593,p11594,p11595,p11596,p11597,p11598,p11599,p11600,p11601,p11602,p11603,p11604,p11605,p11606,p11607,p11608,p11609,p11610,p11611,p11612,p11613,p11614,p11615,p11616,p11617,p11618,p11619,p11620,p11621,p11622,p11623,p11624,p11625,p11626,p11627,p11628,p11629,p11630,p11631,p11632,p11633,p11634,p11635,p11636,p11637,p11638,p11639,p11640,p11641,p11642,p11643,p11644,p11645,p11646,p11647,p11648,p11649,p11650,p11651,p11652,p11653,p11654,p11655,p11656,p11657,p11658,p11659,p11660,p11661,p11662,p11663,p11664,p11665,p11666,p11667,p11668,p11669,p11670,p11671,p11672,p11673,p11674,p11675,p11676,p11677,p11678,p11679,p11680,p11681,p11682,p11683,p11684,p11685,p11686,p11687,p11688,p11689,p11690,p11691,p11692,p11693,p11694,p11695,p11696,p11697,p11698,p11699,p11700,p11701,p11702,p11703,p11704,p11705,p11706,p11707,p11708,p11709,p11710,p11711,p11712,p11713,p11714,p11715,p11716,p11717,p11718,p11719,p11720,p11721,p11722,p11723,p11724,p11725,p11726,p11727,p11728,p11729,p11730,p11731,p11732,p11733,p11734,p11735,p11736,p11737,p11738,p11739,p11740,p11741,p11742,p11743,p11744,p11745,p11746,p11747,p11748,p11749,p11750,p11751,p11752,p11753,p11754,p11755,p11756,p11757,p11758,p11759,p11760,p11761,p11762,p11763,p11764,p11765,p11766,p11767,p11768,p11769,p11770,p11771,p11772,p11773,p11774,p11775,p11776,p11777,p11778,p11779,p11780,p11781,p11782,p11783,p11784,p11785,p11786,p11787,p11788,p11789,p11790,p11791,p11792,p11793,p11794,p11795,p11796,p11797,p11798,p11799,p11800,p11801,p11802,p11803,p11804,p11805,p11806,p11807,p11808,p11809,p11810,p11811,p11812,p11813,p11814,p11815,p11816,p11817,p11818,p11819,p11820,p11821,p11822,p11823,p11824,p11825,p11826,p11827,p11828,p11829,p11830,p11831,p11832,p11833,p11834,p11835,p11836,p11837,p11838,p11839,p11840,p11841,p11842,p11843,p11844,p11845,p11846,p11847,p11848,p11849,p11850,p11851,p11852,p11853,p11854,p11855,p11856,p11857,p11858,p11859,p11860,p11861,p11862,p11863,p11864,p11865,p11866,p11867,p11868,p11869,p11870,p11871,p11872,p11873,p11874,p11875,p11876,p11877,p11878,p11879,p11880,p11881,p11882,p11883,p11884,p11885,p11886,p11887,p11888,p11889,p11890,p11891,p11892,p11893,p11894,p11895,p11896,p11897,p11898,p11899,p11900,p11901,p11902,p11903,p11904,p11905,p11906,p11907,p11908,p11909,p11910,p11911,p11912,p11913,p11914,p11915,p11916,p11917,p11918,p11919,p11920,p11921,p11922,p11923,p11924,p11925,p11926,p11927,p11928,p11929,p11930,p11931,p11932,p11933,p11934,p11935,p11936,p11937,p11938,p11939,p11940,p11941,p11942,p11943,p11944,p11945,p11946,p11947,p11948,p11949,p11950,p11951,p11952,p11953,p11954,p11955,p11956,p11957,p11958,p11959,p11960,p11961,p11962,p11963,p11964,p11965,p11966,p11967,p11968,p11969,p11970,p11971,p11972,p11973,p11974,p11975,p11976,p11977,p11978,p11979,p11980,p11981,p11982,p11983,p11984,p11985,p11986,p11987,p11988,p11989,p11990,p11991,p11992,p11993,p11994,p11995,p11996,p11997,p11998,p11999,p12000,p12001,p12002,p12003,p12004,p12005,p12006,p12007,p12008,p12009,p12010,p12011,p12012,p12013,p12014,p12015,p12016,p12017,p12018,p12019,p12020,p12021,p12022,p12023,p12024,p12025,p12026,p12027,p12028,p12029,p12030,p12031,p12032,p12033,p12034,p12035,p12036,p12037,p12038,p12039,p12040,p12041,p12042,p12043,p12044,p12045,p12046,p12047,p12048,p12049,p12050,p12051,p12052,p12053,p12054,p12055,p12056,p12057,p12058,p12059,p12060,p12061,p12062,p12063,p12064,p12065,p12066,p12067,p12068,p12069,p12070,p12071,p12072,p12073,p12074,p12075,p12076,p12077,p12078,p12079,p12080,p12081,p12082,p12083,p12084,p12085,p12086,p12087,p12088,p12089,p12090,p12091,p12092,p12093,p12094,p12095,p12096,p12097,p12098,p12099,p12100,p12101,p12102,p12103,p12104,p12105,p12106,p12107,p12108,p12109,p12110,p12111,p12112,p12113,p12114,p12115,p12116,p12117,p12118,p12119,p12120,p12121,p12122,p12123,p12124,p12125,p12126,p12127,p12128,p12129,p12130,p12131,p12132,p12133,p12134,p12135,p12136,p12137,p12138,p12139,p12140,p12141,p12142,p12143,p12144,p12145,p12146,p12147,p12148,p12149,p12150,p12151,p12152,p12153,p12154,p12155,p12156,p12157,p12158,p12159,p12160,p12161,p12162,p12163,p12164,p12165,p12166,p12167,p12168,p12169,p12170,p12171,p12172,p12173,p12174,p12175,p12176,p12177,p12178,p12179,p12180,p12181,p12182,p12183,p12184,p12185,p12186,p12187,p12188,p12189,p12190,p12191,p12192,p12193;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_0_8,x[0],y[8]);
and and9(ip_0_9,x[0],y[9]);
and and10(ip_0_10,x[0],y[10]);
and and11(ip_0_11,x[0],y[11]);
and and12(ip_0_12,x[0],y[12]);
and and13(ip_0_13,x[0],y[13]);
and and14(ip_0_14,x[0],y[14]);
and and15(ip_0_15,x[0],y[15]);
and and16(ip_0_16,x[0],y[16]);
and and17(ip_0_17,x[0],y[17]);
and and18(ip_0_18,x[0],y[18]);
and and19(ip_0_19,x[0],y[19]);
and and20(ip_0_20,x[0],y[20]);
and and21(ip_0_21,x[0],y[21]);
and and22(ip_0_22,x[0],y[22]);
and and23(ip_0_23,x[0],y[23]);
and and24(ip_0_24,x[0],y[24]);
and and25(ip_0_25,x[0],y[25]);
and and26(ip_0_26,x[0],y[26]);
and and27(ip_0_27,x[0],y[27]);
and and28(ip_0_28,x[0],y[28]);
and and29(ip_0_29,x[0],y[29]);
and and30(ip_0_30,x[0],y[30]);
and and31(ip_0_31,x[0],y[31]);
and and32(ip_0_32,x[0],y[32]);
and and33(ip_0_33,x[0],y[33]);
and and34(ip_0_34,x[0],y[34]);
and and35(ip_0_35,x[0],y[35]);
and and36(ip_0_36,x[0],y[36]);
and and37(ip_0_37,x[0],y[37]);
and and38(ip_0_38,x[0],y[38]);
and and39(ip_0_39,x[0],y[39]);
and and40(ip_0_40,x[0],y[40]);
and and41(ip_0_41,x[0],y[41]);
and and42(ip_0_42,x[0],y[42]);
and and43(ip_0_43,x[0],y[43]);
and and44(ip_0_44,x[0],y[44]);
and and45(ip_0_45,x[0],y[45]);
and and46(ip_0_46,x[0],y[46]);
and and47(ip_0_47,x[0],y[47]);
and and48(ip_0_48,x[0],y[48]);
and and49(ip_0_49,x[0],y[49]);
and and50(ip_0_50,x[0],y[50]);
and and51(ip_0_51,x[0],y[51]);
and and52(ip_0_52,x[0],y[52]);
and and53(ip_0_53,x[0],y[53]);
and and54(ip_0_54,x[0],y[54]);
and and55(ip_0_55,x[0],y[55]);
and and56(ip_0_56,x[0],y[56]);
and and57(ip_0_57,x[0],y[57]);
and and58(ip_0_58,x[0],y[58]);
and and59(ip_0_59,x[0],y[59]);
and and60(ip_0_60,x[0],y[60]);
and and61(ip_0_61,x[0],y[61]);
and and62(ip_0_62,x[0],y[62]);
and and63(ip_0_63,x[0],y[63]);
and and64(ip_1_0,x[1],y[0]);
and and65(ip_1_1,x[1],y[1]);
and and66(ip_1_2,x[1],y[2]);
and and67(ip_1_3,x[1],y[3]);
and and68(ip_1_4,x[1],y[4]);
and and69(ip_1_5,x[1],y[5]);
and and70(ip_1_6,x[1],y[6]);
and and71(ip_1_7,x[1],y[7]);
and and72(ip_1_8,x[1],y[8]);
and and73(ip_1_9,x[1],y[9]);
and and74(ip_1_10,x[1],y[10]);
and and75(ip_1_11,x[1],y[11]);
and and76(ip_1_12,x[1],y[12]);
and and77(ip_1_13,x[1],y[13]);
and and78(ip_1_14,x[1],y[14]);
and and79(ip_1_15,x[1],y[15]);
and and80(ip_1_16,x[1],y[16]);
and and81(ip_1_17,x[1],y[17]);
and and82(ip_1_18,x[1],y[18]);
and and83(ip_1_19,x[1],y[19]);
and and84(ip_1_20,x[1],y[20]);
and and85(ip_1_21,x[1],y[21]);
and and86(ip_1_22,x[1],y[22]);
and and87(ip_1_23,x[1],y[23]);
and and88(ip_1_24,x[1],y[24]);
and and89(ip_1_25,x[1],y[25]);
and and90(ip_1_26,x[1],y[26]);
and and91(ip_1_27,x[1],y[27]);
and and92(ip_1_28,x[1],y[28]);
and and93(ip_1_29,x[1],y[29]);
and and94(ip_1_30,x[1],y[30]);
and and95(ip_1_31,x[1],y[31]);
and and96(ip_1_32,x[1],y[32]);
and and97(ip_1_33,x[1],y[33]);
and and98(ip_1_34,x[1],y[34]);
and and99(ip_1_35,x[1],y[35]);
and and100(ip_1_36,x[1],y[36]);
and and101(ip_1_37,x[1],y[37]);
and and102(ip_1_38,x[1],y[38]);
and and103(ip_1_39,x[1],y[39]);
and and104(ip_1_40,x[1],y[40]);
and and105(ip_1_41,x[1],y[41]);
and and106(ip_1_42,x[1],y[42]);
and and107(ip_1_43,x[1],y[43]);
and and108(ip_1_44,x[1],y[44]);
and and109(ip_1_45,x[1],y[45]);
and and110(ip_1_46,x[1],y[46]);
and and111(ip_1_47,x[1],y[47]);
and and112(ip_1_48,x[1],y[48]);
and and113(ip_1_49,x[1],y[49]);
and and114(ip_1_50,x[1],y[50]);
and and115(ip_1_51,x[1],y[51]);
and and116(ip_1_52,x[1],y[52]);
and and117(ip_1_53,x[1],y[53]);
and and118(ip_1_54,x[1],y[54]);
and and119(ip_1_55,x[1],y[55]);
and and120(ip_1_56,x[1],y[56]);
and and121(ip_1_57,x[1],y[57]);
and and122(ip_1_58,x[1],y[58]);
and and123(ip_1_59,x[1],y[59]);
and and124(ip_1_60,x[1],y[60]);
and and125(ip_1_61,x[1],y[61]);
and and126(ip_1_62,x[1],y[62]);
and and127(ip_1_63,x[1],y[63]);
and and128(ip_2_0,x[2],y[0]);
and and129(ip_2_1,x[2],y[1]);
and and130(ip_2_2,x[2],y[2]);
and and131(ip_2_3,x[2],y[3]);
and and132(ip_2_4,x[2],y[4]);
and and133(ip_2_5,x[2],y[5]);
and and134(ip_2_6,x[2],y[6]);
and and135(ip_2_7,x[2],y[7]);
and and136(ip_2_8,x[2],y[8]);
and and137(ip_2_9,x[2],y[9]);
and and138(ip_2_10,x[2],y[10]);
and and139(ip_2_11,x[2],y[11]);
and and140(ip_2_12,x[2],y[12]);
and and141(ip_2_13,x[2],y[13]);
and and142(ip_2_14,x[2],y[14]);
and and143(ip_2_15,x[2],y[15]);
and and144(ip_2_16,x[2],y[16]);
and and145(ip_2_17,x[2],y[17]);
and and146(ip_2_18,x[2],y[18]);
and and147(ip_2_19,x[2],y[19]);
and and148(ip_2_20,x[2],y[20]);
and and149(ip_2_21,x[2],y[21]);
and and150(ip_2_22,x[2],y[22]);
and and151(ip_2_23,x[2],y[23]);
and and152(ip_2_24,x[2],y[24]);
and and153(ip_2_25,x[2],y[25]);
and and154(ip_2_26,x[2],y[26]);
and and155(ip_2_27,x[2],y[27]);
and and156(ip_2_28,x[2],y[28]);
and and157(ip_2_29,x[2],y[29]);
and and158(ip_2_30,x[2],y[30]);
and and159(ip_2_31,x[2],y[31]);
and and160(ip_2_32,x[2],y[32]);
and and161(ip_2_33,x[2],y[33]);
and and162(ip_2_34,x[2],y[34]);
and and163(ip_2_35,x[2],y[35]);
and and164(ip_2_36,x[2],y[36]);
and and165(ip_2_37,x[2],y[37]);
and and166(ip_2_38,x[2],y[38]);
and and167(ip_2_39,x[2],y[39]);
and and168(ip_2_40,x[2],y[40]);
and and169(ip_2_41,x[2],y[41]);
and and170(ip_2_42,x[2],y[42]);
and and171(ip_2_43,x[2],y[43]);
and and172(ip_2_44,x[2],y[44]);
and and173(ip_2_45,x[2],y[45]);
and and174(ip_2_46,x[2],y[46]);
and and175(ip_2_47,x[2],y[47]);
and and176(ip_2_48,x[2],y[48]);
and and177(ip_2_49,x[2],y[49]);
and and178(ip_2_50,x[2],y[50]);
and and179(ip_2_51,x[2],y[51]);
and and180(ip_2_52,x[2],y[52]);
and and181(ip_2_53,x[2],y[53]);
and and182(ip_2_54,x[2],y[54]);
and and183(ip_2_55,x[2],y[55]);
and and184(ip_2_56,x[2],y[56]);
and and185(ip_2_57,x[2],y[57]);
and and186(ip_2_58,x[2],y[58]);
and and187(ip_2_59,x[2],y[59]);
and and188(ip_2_60,x[2],y[60]);
and and189(ip_2_61,x[2],y[61]);
and and190(ip_2_62,x[2],y[62]);
and and191(ip_2_63,x[2],y[63]);
and and192(ip_3_0,x[3],y[0]);
and and193(ip_3_1,x[3],y[1]);
and and194(ip_3_2,x[3],y[2]);
and and195(ip_3_3,x[3],y[3]);
and and196(ip_3_4,x[3],y[4]);
and and197(ip_3_5,x[3],y[5]);
and and198(ip_3_6,x[3],y[6]);
and and199(ip_3_7,x[3],y[7]);
and and200(ip_3_8,x[3],y[8]);
and and201(ip_3_9,x[3],y[9]);
and and202(ip_3_10,x[3],y[10]);
and and203(ip_3_11,x[3],y[11]);
and and204(ip_3_12,x[3],y[12]);
and and205(ip_3_13,x[3],y[13]);
and and206(ip_3_14,x[3],y[14]);
and and207(ip_3_15,x[3],y[15]);
and and208(ip_3_16,x[3],y[16]);
and and209(ip_3_17,x[3],y[17]);
and and210(ip_3_18,x[3],y[18]);
and and211(ip_3_19,x[3],y[19]);
and and212(ip_3_20,x[3],y[20]);
and and213(ip_3_21,x[3],y[21]);
and and214(ip_3_22,x[3],y[22]);
and and215(ip_3_23,x[3],y[23]);
and and216(ip_3_24,x[3],y[24]);
and and217(ip_3_25,x[3],y[25]);
and and218(ip_3_26,x[3],y[26]);
and and219(ip_3_27,x[3],y[27]);
and and220(ip_3_28,x[3],y[28]);
and and221(ip_3_29,x[3],y[29]);
and and222(ip_3_30,x[3],y[30]);
and and223(ip_3_31,x[3],y[31]);
and and224(ip_3_32,x[3],y[32]);
and and225(ip_3_33,x[3],y[33]);
and and226(ip_3_34,x[3],y[34]);
and and227(ip_3_35,x[3],y[35]);
and and228(ip_3_36,x[3],y[36]);
and and229(ip_3_37,x[3],y[37]);
and and230(ip_3_38,x[3],y[38]);
and and231(ip_3_39,x[3],y[39]);
and and232(ip_3_40,x[3],y[40]);
and and233(ip_3_41,x[3],y[41]);
and and234(ip_3_42,x[3],y[42]);
and and235(ip_3_43,x[3],y[43]);
and and236(ip_3_44,x[3],y[44]);
and and237(ip_3_45,x[3],y[45]);
and and238(ip_3_46,x[3],y[46]);
and and239(ip_3_47,x[3],y[47]);
and and240(ip_3_48,x[3],y[48]);
and and241(ip_3_49,x[3],y[49]);
and and242(ip_3_50,x[3],y[50]);
and and243(ip_3_51,x[3],y[51]);
and and244(ip_3_52,x[3],y[52]);
and and245(ip_3_53,x[3],y[53]);
and and246(ip_3_54,x[3],y[54]);
and and247(ip_3_55,x[3],y[55]);
and and248(ip_3_56,x[3],y[56]);
and and249(ip_3_57,x[3],y[57]);
and and250(ip_3_58,x[3],y[58]);
and and251(ip_3_59,x[3],y[59]);
and and252(ip_3_60,x[3],y[60]);
and and253(ip_3_61,x[3],y[61]);
and and254(ip_3_62,x[3],y[62]);
and and255(ip_3_63,x[3],y[63]);
and and256(ip_4_0,x[4],y[0]);
and and257(ip_4_1,x[4],y[1]);
and and258(ip_4_2,x[4],y[2]);
and and259(ip_4_3,x[4],y[3]);
and and260(ip_4_4,x[4],y[4]);
and and261(ip_4_5,x[4],y[5]);
and and262(ip_4_6,x[4],y[6]);
and and263(ip_4_7,x[4],y[7]);
and and264(ip_4_8,x[4],y[8]);
and and265(ip_4_9,x[4],y[9]);
and and266(ip_4_10,x[4],y[10]);
and and267(ip_4_11,x[4],y[11]);
and and268(ip_4_12,x[4],y[12]);
and and269(ip_4_13,x[4],y[13]);
and and270(ip_4_14,x[4],y[14]);
and and271(ip_4_15,x[4],y[15]);
and and272(ip_4_16,x[4],y[16]);
and and273(ip_4_17,x[4],y[17]);
and and274(ip_4_18,x[4],y[18]);
and and275(ip_4_19,x[4],y[19]);
and and276(ip_4_20,x[4],y[20]);
and and277(ip_4_21,x[4],y[21]);
and and278(ip_4_22,x[4],y[22]);
and and279(ip_4_23,x[4],y[23]);
and and280(ip_4_24,x[4],y[24]);
and and281(ip_4_25,x[4],y[25]);
and and282(ip_4_26,x[4],y[26]);
and and283(ip_4_27,x[4],y[27]);
and and284(ip_4_28,x[4],y[28]);
and and285(ip_4_29,x[4],y[29]);
and and286(ip_4_30,x[4],y[30]);
and and287(ip_4_31,x[4],y[31]);
and and288(ip_4_32,x[4],y[32]);
and and289(ip_4_33,x[4],y[33]);
and and290(ip_4_34,x[4],y[34]);
and and291(ip_4_35,x[4],y[35]);
and and292(ip_4_36,x[4],y[36]);
and and293(ip_4_37,x[4],y[37]);
and and294(ip_4_38,x[4],y[38]);
and and295(ip_4_39,x[4],y[39]);
and and296(ip_4_40,x[4],y[40]);
and and297(ip_4_41,x[4],y[41]);
and and298(ip_4_42,x[4],y[42]);
and and299(ip_4_43,x[4],y[43]);
and and300(ip_4_44,x[4],y[44]);
and and301(ip_4_45,x[4],y[45]);
and and302(ip_4_46,x[4],y[46]);
and and303(ip_4_47,x[4],y[47]);
and and304(ip_4_48,x[4],y[48]);
and and305(ip_4_49,x[4],y[49]);
and and306(ip_4_50,x[4],y[50]);
and and307(ip_4_51,x[4],y[51]);
and and308(ip_4_52,x[4],y[52]);
and and309(ip_4_53,x[4],y[53]);
and and310(ip_4_54,x[4],y[54]);
and and311(ip_4_55,x[4],y[55]);
and and312(ip_4_56,x[4],y[56]);
and and313(ip_4_57,x[4],y[57]);
and and314(ip_4_58,x[4],y[58]);
and and315(ip_4_59,x[4],y[59]);
and and316(ip_4_60,x[4],y[60]);
and and317(ip_4_61,x[4],y[61]);
and and318(ip_4_62,x[4],y[62]);
and and319(ip_4_63,x[4],y[63]);
and and320(ip_5_0,x[5],y[0]);
and and321(ip_5_1,x[5],y[1]);
and and322(ip_5_2,x[5],y[2]);
and and323(ip_5_3,x[5],y[3]);
and and324(ip_5_4,x[5],y[4]);
and and325(ip_5_5,x[5],y[5]);
and and326(ip_5_6,x[5],y[6]);
and and327(ip_5_7,x[5],y[7]);
and and328(ip_5_8,x[5],y[8]);
and and329(ip_5_9,x[5],y[9]);
and and330(ip_5_10,x[5],y[10]);
and and331(ip_5_11,x[5],y[11]);
and and332(ip_5_12,x[5],y[12]);
and and333(ip_5_13,x[5],y[13]);
and and334(ip_5_14,x[5],y[14]);
and and335(ip_5_15,x[5],y[15]);
and and336(ip_5_16,x[5],y[16]);
and and337(ip_5_17,x[5],y[17]);
and and338(ip_5_18,x[5],y[18]);
and and339(ip_5_19,x[5],y[19]);
and and340(ip_5_20,x[5],y[20]);
and and341(ip_5_21,x[5],y[21]);
and and342(ip_5_22,x[5],y[22]);
and and343(ip_5_23,x[5],y[23]);
and and344(ip_5_24,x[5],y[24]);
and and345(ip_5_25,x[5],y[25]);
and and346(ip_5_26,x[5],y[26]);
and and347(ip_5_27,x[5],y[27]);
and and348(ip_5_28,x[5],y[28]);
and and349(ip_5_29,x[5],y[29]);
and and350(ip_5_30,x[5],y[30]);
and and351(ip_5_31,x[5],y[31]);
and and352(ip_5_32,x[5],y[32]);
and and353(ip_5_33,x[5],y[33]);
and and354(ip_5_34,x[5],y[34]);
and and355(ip_5_35,x[5],y[35]);
and and356(ip_5_36,x[5],y[36]);
and and357(ip_5_37,x[5],y[37]);
and and358(ip_5_38,x[5],y[38]);
and and359(ip_5_39,x[5],y[39]);
and and360(ip_5_40,x[5],y[40]);
and and361(ip_5_41,x[5],y[41]);
and and362(ip_5_42,x[5],y[42]);
and and363(ip_5_43,x[5],y[43]);
and and364(ip_5_44,x[5],y[44]);
and and365(ip_5_45,x[5],y[45]);
and and366(ip_5_46,x[5],y[46]);
and and367(ip_5_47,x[5],y[47]);
and and368(ip_5_48,x[5],y[48]);
and and369(ip_5_49,x[5],y[49]);
and and370(ip_5_50,x[5],y[50]);
and and371(ip_5_51,x[5],y[51]);
and and372(ip_5_52,x[5],y[52]);
and and373(ip_5_53,x[5],y[53]);
and and374(ip_5_54,x[5],y[54]);
and and375(ip_5_55,x[5],y[55]);
and and376(ip_5_56,x[5],y[56]);
and and377(ip_5_57,x[5],y[57]);
and and378(ip_5_58,x[5],y[58]);
and and379(ip_5_59,x[5],y[59]);
and and380(ip_5_60,x[5],y[60]);
and and381(ip_5_61,x[5],y[61]);
and and382(ip_5_62,x[5],y[62]);
and and383(ip_5_63,x[5],y[63]);
and and384(ip_6_0,x[6],y[0]);
and and385(ip_6_1,x[6],y[1]);
and and386(ip_6_2,x[6],y[2]);
and and387(ip_6_3,x[6],y[3]);
and and388(ip_6_4,x[6],y[4]);
and and389(ip_6_5,x[6],y[5]);
and and390(ip_6_6,x[6],y[6]);
and and391(ip_6_7,x[6],y[7]);
and and392(ip_6_8,x[6],y[8]);
and and393(ip_6_9,x[6],y[9]);
and and394(ip_6_10,x[6],y[10]);
and and395(ip_6_11,x[6],y[11]);
and and396(ip_6_12,x[6],y[12]);
and and397(ip_6_13,x[6],y[13]);
and and398(ip_6_14,x[6],y[14]);
and and399(ip_6_15,x[6],y[15]);
and and400(ip_6_16,x[6],y[16]);
and and401(ip_6_17,x[6],y[17]);
and and402(ip_6_18,x[6],y[18]);
and and403(ip_6_19,x[6],y[19]);
and and404(ip_6_20,x[6],y[20]);
and and405(ip_6_21,x[6],y[21]);
and and406(ip_6_22,x[6],y[22]);
and and407(ip_6_23,x[6],y[23]);
and and408(ip_6_24,x[6],y[24]);
and and409(ip_6_25,x[6],y[25]);
and and410(ip_6_26,x[6],y[26]);
and and411(ip_6_27,x[6],y[27]);
and and412(ip_6_28,x[6],y[28]);
and and413(ip_6_29,x[6],y[29]);
and and414(ip_6_30,x[6],y[30]);
and and415(ip_6_31,x[6],y[31]);
and and416(ip_6_32,x[6],y[32]);
and and417(ip_6_33,x[6],y[33]);
and and418(ip_6_34,x[6],y[34]);
and and419(ip_6_35,x[6],y[35]);
and and420(ip_6_36,x[6],y[36]);
and and421(ip_6_37,x[6],y[37]);
and and422(ip_6_38,x[6],y[38]);
and and423(ip_6_39,x[6],y[39]);
and and424(ip_6_40,x[6],y[40]);
and and425(ip_6_41,x[6],y[41]);
and and426(ip_6_42,x[6],y[42]);
and and427(ip_6_43,x[6],y[43]);
and and428(ip_6_44,x[6],y[44]);
and and429(ip_6_45,x[6],y[45]);
and and430(ip_6_46,x[6],y[46]);
and and431(ip_6_47,x[6],y[47]);
and and432(ip_6_48,x[6],y[48]);
and and433(ip_6_49,x[6],y[49]);
and and434(ip_6_50,x[6],y[50]);
and and435(ip_6_51,x[6],y[51]);
and and436(ip_6_52,x[6],y[52]);
and and437(ip_6_53,x[6],y[53]);
and and438(ip_6_54,x[6],y[54]);
and and439(ip_6_55,x[6],y[55]);
and and440(ip_6_56,x[6],y[56]);
and and441(ip_6_57,x[6],y[57]);
and and442(ip_6_58,x[6],y[58]);
and and443(ip_6_59,x[6],y[59]);
and and444(ip_6_60,x[6],y[60]);
and and445(ip_6_61,x[6],y[61]);
and and446(ip_6_62,x[6],y[62]);
and and447(ip_6_63,x[6],y[63]);
and and448(ip_7_0,x[7],y[0]);
and and449(ip_7_1,x[7],y[1]);
and and450(ip_7_2,x[7],y[2]);
and and451(ip_7_3,x[7],y[3]);
and and452(ip_7_4,x[7],y[4]);
and and453(ip_7_5,x[7],y[5]);
and and454(ip_7_6,x[7],y[6]);
and and455(ip_7_7,x[7],y[7]);
and and456(ip_7_8,x[7],y[8]);
and and457(ip_7_9,x[7],y[9]);
and and458(ip_7_10,x[7],y[10]);
and and459(ip_7_11,x[7],y[11]);
and and460(ip_7_12,x[7],y[12]);
and and461(ip_7_13,x[7],y[13]);
and and462(ip_7_14,x[7],y[14]);
and and463(ip_7_15,x[7],y[15]);
and and464(ip_7_16,x[7],y[16]);
and and465(ip_7_17,x[7],y[17]);
and and466(ip_7_18,x[7],y[18]);
and and467(ip_7_19,x[7],y[19]);
and and468(ip_7_20,x[7],y[20]);
and and469(ip_7_21,x[7],y[21]);
and and470(ip_7_22,x[7],y[22]);
and and471(ip_7_23,x[7],y[23]);
and and472(ip_7_24,x[7],y[24]);
and and473(ip_7_25,x[7],y[25]);
and and474(ip_7_26,x[7],y[26]);
and and475(ip_7_27,x[7],y[27]);
and and476(ip_7_28,x[7],y[28]);
and and477(ip_7_29,x[7],y[29]);
and and478(ip_7_30,x[7],y[30]);
and and479(ip_7_31,x[7],y[31]);
and and480(ip_7_32,x[7],y[32]);
and and481(ip_7_33,x[7],y[33]);
and and482(ip_7_34,x[7],y[34]);
and and483(ip_7_35,x[7],y[35]);
and and484(ip_7_36,x[7],y[36]);
and and485(ip_7_37,x[7],y[37]);
and and486(ip_7_38,x[7],y[38]);
and and487(ip_7_39,x[7],y[39]);
and and488(ip_7_40,x[7],y[40]);
and and489(ip_7_41,x[7],y[41]);
and and490(ip_7_42,x[7],y[42]);
and and491(ip_7_43,x[7],y[43]);
and and492(ip_7_44,x[7],y[44]);
and and493(ip_7_45,x[7],y[45]);
and and494(ip_7_46,x[7],y[46]);
and and495(ip_7_47,x[7],y[47]);
and and496(ip_7_48,x[7],y[48]);
and and497(ip_7_49,x[7],y[49]);
and and498(ip_7_50,x[7],y[50]);
and and499(ip_7_51,x[7],y[51]);
and and500(ip_7_52,x[7],y[52]);
and and501(ip_7_53,x[7],y[53]);
and and502(ip_7_54,x[7],y[54]);
and and503(ip_7_55,x[7],y[55]);
and and504(ip_7_56,x[7],y[56]);
and and505(ip_7_57,x[7],y[57]);
and and506(ip_7_58,x[7],y[58]);
and and507(ip_7_59,x[7],y[59]);
and and508(ip_7_60,x[7],y[60]);
and and509(ip_7_61,x[7],y[61]);
and and510(ip_7_62,x[7],y[62]);
and and511(ip_7_63,x[7],y[63]);
and and512(ip_8_0,x[8],y[0]);
and and513(ip_8_1,x[8],y[1]);
and and514(ip_8_2,x[8],y[2]);
and and515(ip_8_3,x[8],y[3]);
and and516(ip_8_4,x[8],y[4]);
and and517(ip_8_5,x[8],y[5]);
and and518(ip_8_6,x[8],y[6]);
and and519(ip_8_7,x[8],y[7]);
and and520(ip_8_8,x[8],y[8]);
and and521(ip_8_9,x[8],y[9]);
and and522(ip_8_10,x[8],y[10]);
and and523(ip_8_11,x[8],y[11]);
and and524(ip_8_12,x[8],y[12]);
and and525(ip_8_13,x[8],y[13]);
and and526(ip_8_14,x[8],y[14]);
and and527(ip_8_15,x[8],y[15]);
and and528(ip_8_16,x[8],y[16]);
and and529(ip_8_17,x[8],y[17]);
and and530(ip_8_18,x[8],y[18]);
and and531(ip_8_19,x[8],y[19]);
and and532(ip_8_20,x[8],y[20]);
and and533(ip_8_21,x[8],y[21]);
and and534(ip_8_22,x[8],y[22]);
and and535(ip_8_23,x[8],y[23]);
and and536(ip_8_24,x[8],y[24]);
and and537(ip_8_25,x[8],y[25]);
and and538(ip_8_26,x[8],y[26]);
and and539(ip_8_27,x[8],y[27]);
and and540(ip_8_28,x[8],y[28]);
and and541(ip_8_29,x[8],y[29]);
and and542(ip_8_30,x[8],y[30]);
and and543(ip_8_31,x[8],y[31]);
and and544(ip_8_32,x[8],y[32]);
and and545(ip_8_33,x[8],y[33]);
and and546(ip_8_34,x[8],y[34]);
and and547(ip_8_35,x[8],y[35]);
and and548(ip_8_36,x[8],y[36]);
and and549(ip_8_37,x[8],y[37]);
and and550(ip_8_38,x[8],y[38]);
and and551(ip_8_39,x[8],y[39]);
and and552(ip_8_40,x[8],y[40]);
and and553(ip_8_41,x[8],y[41]);
and and554(ip_8_42,x[8],y[42]);
and and555(ip_8_43,x[8],y[43]);
and and556(ip_8_44,x[8],y[44]);
and and557(ip_8_45,x[8],y[45]);
and and558(ip_8_46,x[8],y[46]);
and and559(ip_8_47,x[8],y[47]);
and and560(ip_8_48,x[8],y[48]);
and and561(ip_8_49,x[8],y[49]);
and and562(ip_8_50,x[8],y[50]);
and and563(ip_8_51,x[8],y[51]);
and and564(ip_8_52,x[8],y[52]);
and and565(ip_8_53,x[8],y[53]);
and and566(ip_8_54,x[8],y[54]);
and and567(ip_8_55,x[8],y[55]);
and and568(ip_8_56,x[8],y[56]);
and and569(ip_8_57,x[8],y[57]);
and and570(ip_8_58,x[8],y[58]);
and and571(ip_8_59,x[8],y[59]);
and and572(ip_8_60,x[8],y[60]);
and and573(ip_8_61,x[8],y[61]);
and and574(ip_8_62,x[8],y[62]);
and and575(ip_8_63,x[8],y[63]);
and and576(ip_9_0,x[9],y[0]);
and and577(ip_9_1,x[9],y[1]);
and and578(ip_9_2,x[9],y[2]);
and and579(ip_9_3,x[9],y[3]);
and and580(ip_9_4,x[9],y[4]);
and and581(ip_9_5,x[9],y[5]);
and and582(ip_9_6,x[9],y[6]);
and and583(ip_9_7,x[9],y[7]);
and and584(ip_9_8,x[9],y[8]);
and and585(ip_9_9,x[9],y[9]);
and and586(ip_9_10,x[9],y[10]);
and and587(ip_9_11,x[9],y[11]);
and and588(ip_9_12,x[9],y[12]);
and and589(ip_9_13,x[9],y[13]);
and and590(ip_9_14,x[9],y[14]);
and and591(ip_9_15,x[9],y[15]);
and and592(ip_9_16,x[9],y[16]);
and and593(ip_9_17,x[9],y[17]);
and and594(ip_9_18,x[9],y[18]);
and and595(ip_9_19,x[9],y[19]);
and and596(ip_9_20,x[9],y[20]);
and and597(ip_9_21,x[9],y[21]);
and and598(ip_9_22,x[9],y[22]);
and and599(ip_9_23,x[9],y[23]);
and and600(ip_9_24,x[9],y[24]);
and and601(ip_9_25,x[9],y[25]);
and and602(ip_9_26,x[9],y[26]);
and and603(ip_9_27,x[9],y[27]);
and and604(ip_9_28,x[9],y[28]);
and and605(ip_9_29,x[9],y[29]);
and and606(ip_9_30,x[9],y[30]);
and and607(ip_9_31,x[9],y[31]);
and and608(ip_9_32,x[9],y[32]);
and and609(ip_9_33,x[9],y[33]);
and and610(ip_9_34,x[9],y[34]);
and and611(ip_9_35,x[9],y[35]);
and and612(ip_9_36,x[9],y[36]);
and and613(ip_9_37,x[9],y[37]);
and and614(ip_9_38,x[9],y[38]);
and and615(ip_9_39,x[9],y[39]);
and and616(ip_9_40,x[9],y[40]);
and and617(ip_9_41,x[9],y[41]);
and and618(ip_9_42,x[9],y[42]);
and and619(ip_9_43,x[9],y[43]);
and and620(ip_9_44,x[9],y[44]);
and and621(ip_9_45,x[9],y[45]);
and and622(ip_9_46,x[9],y[46]);
and and623(ip_9_47,x[9],y[47]);
and and624(ip_9_48,x[9],y[48]);
and and625(ip_9_49,x[9],y[49]);
and and626(ip_9_50,x[9],y[50]);
and and627(ip_9_51,x[9],y[51]);
and and628(ip_9_52,x[9],y[52]);
and and629(ip_9_53,x[9],y[53]);
and and630(ip_9_54,x[9],y[54]);
and and631(ip_9_55,x[9],y[55]);
and and632(ip_9_56,x[9],y[56]);
and and633(ip_9_57,x[9],y[57]);
and and634(ip_9_58,x[9],y[58]);
and and635(ip_9_59,x[9],y[59]);
and and636(ip_9_60,x[9],y[60]);
and and637(ip_9_61,x[9],y[61]);
and and638(ip_9_62,x[9],y[62]);
and and639(ip_9_63,x[9],y[63]);
and and640(ip_10_0,x[10],y[0]);
and and641(ip_10_1,x[10],y[1]);
and and642(ip_10_2,x[10],y[2]);
and and643(ip_10_3,x[10],y[3]);
and and644(ip_10_4,x[10],y[4]);
and and645(ip_10_5,x[10],y[5]);
and and646(ip_10_6,x[10],y[6]);
and and647(ip_10_7,x[10],y[7]);
and and648(ip_10_8,x[10],y[8]);
and and649(ip_10_9,x[10],y[9]);
and and650(ip_10_10,x[10],y[10]);
and and651(ip_10_11,x[10],y[11]);
and and652(ip_10_12,x[10],y[12]);
and and653(ip_10_13,x[10],y[13]);
and and654(ip_10_14,x[10],y[14]);
and and655(ip_10_15,x[10],y[15]);
and and656(ip_10_16,x[10],y[16]);
and and657(ip_10_17,x[10],y[17]);
and and658(ip_10_18,x[10],y[18]);
and and659(ip_10_19,x[10],y[19]);
and and660(ip_10_20,x[10],y[20]);
and and661(ip_10_21,x[10],y[21]);
and and662(ip_10_22,x[10],y[22]);
and and663(ip_10_23,x[10],y[23]);
and and664(ip_10_24,x[10],y[24]);
and and665(ip_10_25,x[10],y[25]);
and and666(ip_10_26,x[10],y[26]);
and and667(ip_10_27,x[10],y[27]);
and and668(ip_10_28,x[10],y[28]);
and and669(ip_10_29,x[10],y[29]);
and and670(ip_10_30,x[10],y[30]);
and and671(ip_10_31,x[10],y[31]);
and and672(ip_10_32,x[10],y[32]);
and and673(ip_10_33,x[10],y[33]);
and and674(ip_10_34,x[10],y[34]);
and and675(ip_10_35,x[10],y[35]);
and and676(ip_10_36,x[10],y[36]);
and and677(ip_10_37,x[10],y[37]);
and and678(ip_10_38,x[10],y[38]);
and and679(ip_10_39,x[10],y[39]);
and and680(ip_10_40,x[10],y[40]);
and and681(ip_10_41,x[10],y[41]);
and and682(ip_10_42,x[10],y[42]);
and and683(ip_10_43,x[10],y[43]);
and and684(ip_10_44,x[10],y[44]);
and and685(ip_10_45,x[10],y[45]);
and and686(ip_10_46,x[10],y[46]);
and and687(ip_10_47,x[10],y[47]);
and and688(ip_10_48,x[10],y[48]);
and and689(ip_10_49,x[10],y[49]);
and and690(ip_10_50,x[10],y[50]);
and and691(ip_10_51,x[10],y[51]);
and and692(ip_10_52,x[10],y[52]);
and and693(ip_10_53,x[10],y[53]);
and and694(ip_10_54,x[10],y[54]);
and and695(ip_10_55,x[10],y[55]);
and and696(ip_10_56,x[10],y[56]);
and and697(ip_10_57,x[10],y[57]);
and and698(ip_10_58,x[10],y[58]);
and and699(ip_10_59,x[10],y[59]);
and and700(ip_10_60,x[10],y[60]);
and and701(ip_10_61,x[10],y[61]);
and and702(ip_10_62,x[10],y[62]);
and and703(ip_10_63,x[10],y[63]);
and and704(ip_11_0,x[11],y[0]);
and and705(ip_11_1,x[11],y[1]);
and and706(ip_11_2,x[11],y[2]);
and and707(ip_11_3,x[11],y[3]);
and and708(ip_11_4,x[11],y[4]);
and and709(ip_11_5,x[11],y[5]);
and and710(ip_11_6,x[11],y[6]);
and and711(ip_11_7,x[11],y[7]);
and and712(ip_11_8,x[11],y[8]);
and and713(ip_11_9,x[11],y[9]);
and and714(ip_11_10,x[11],y[10]);
and and715(ip_11_11,x[11],y[11]);
and and716(ip_11_12,x[11],y[12]);
and and717(ip_11_13,x[11],y[13]);
and and718(ip_11_14,x[11],y[14]);
and and719(ip_11_15,x[11],y[15]);
and and720(ip_11_16,x[11],y[16]);
and and721(ip_11_17,x[11],y[17]);
and and722(ip_11_18,x[11],y[18]);
and and723(ip_11_19,x[11],y[19]);
and and724(ip_11_20,x[11],y[20]);
and and725(ip_11_21,x[11],y[21]);
and and726(ip_11_22,x[11],y[22]);
and and727(ip_11_23,x[11],y[23]);
and and728(ip_11_24,x[11],y[24]);
and and729(ip_11_25,x[11],y[25]);
and and730(ip_11_26,x[11],y[26]);
and and731(ip_11_27,x[11],y[27]);
and and732(ip_11_28,x[11],y[28]);
and and733(ip_11_29,x[11],y[29]);
and and734(ip_11_30,x[11],y[30]);
and and735(ip_11_31,x[11],y[31]);
and and736(ip_11_32,x[11],y[32]);
and and737(ip_11_33,x[11],y[33]);
and and738(ip_11_34,x[11],y[34]);
and and739(ip_11_35,x[11],y[35]);
and and740(ip_11_36,x[11],y[36]);
and and741(ip_11_37,x[11],y[37]);
and and742(ip_11_38,x[11],y[38]);
and and743(ip_11_39,x[11],y[39]);
and and744(ip_11_40,x[11],y[40]);
and and745(ip_11_41,x[11],y[41]);
and and746(ip_11_42,x[11],y[42]);
and and747(ip_11_43,x[11],y[43]);
and and748(ip_11_44,x[11],y[44]);
and and749(ip_11_45,x[11],y[45]);
and and750(ip_11_46,x[11],y[46]);
and and751(ip_11_47,x[11],y[47]);
and and752(ip_11_48,x[11],y[48]);
and and753(ip_11_49,x[11],y[49]);
and and754(ip_11_50,x[11],y[50]);
and and755(ip_11_51,x[11],y[51]);
and and756(ip_11_52,x[11],y[52]);
and and757(ip_11_53,x[11],y[53]);
and and758(ip_11_54,x[11],y[54]);
and and759(ip_11_55,x[11],y[55]);
and and760(ip_11_56,x[11],y[56]);
and and761(ip_11_57,x[11],y[57]);
and and762(ip_11_58,x[11],y[58]);
and and763(ip_11_59,x[11],y[59]);
and and764(ip_11_60,x[11],y[60]);
and and765(ip_11_61,x[11],y[61]);
and and766(ip_11_62,x[11],y[62]);
and and767(ip_11_63,x[11],y[63]);
and and768(ip_12_0,x[12],y[0]);
and and769(ip_12_1,x[12],y[1]);
and and770(ip_12_2,x[12],y[2]);
and and771(ip_12_3,x[12],y[3]);
and and772(ip_12_4,x[12],y[4]);
and and773(ip_12_5,x[12],y[5]);
and and774(ip_12_6,x[12],y[6]);
and and775(ip_12_7,x[12],y[7]);
and and776(ip_12_8,x[12],y[8]);
and and777(ip_12_9,x[12],y[9]);
and and778(ip_12_10,x[12],y[10]);
and and779(ip_12_11,x[12],y[11]);
and and780(ip_12_12,x[12],y[12]);
and and781(ip_12_13,x[12],y[13]);
and and782(ip_12_14,x[12],y[14]);
and and783(ip_12_15,x[12],y[15]);
and and784(ip_12_16,x[12],y[16]);
and and785(ip_12_17,x[12],y[17]);
and and786(ip_12_18,x[12],y[18]);
and and787(ip_12_19,x[12],y[19]);
and and788(ip_12_20,x[12],y[20]);
and and789(ip_12_21,x[12],y[21]);
and and790(ip_12_22,x[12],y[22]);
and and791(ip_12_23,x[12],y[23]);
and and792(ip_12_24,x[12],y[24]);
and and793(ip_12_25,x[12],y[25]);
and and794(ip_12_26,x[12],y[26]);
and and795(ip_12_27,x[12],y[27]);
and and796(ip_12_28,x[12],y[28]);
and and797(ip_12_29,x[12],y[29]);
and and798(ip_12_30,x[12],y[30]);
and and799(ip_12_31,x[12],y[31]);
and and800(ip_12_32,x[12],y[32]);
and and801(ip_12_33,x[12],y[33]);
and and802(ip_12_34,x[12],y[34]);
and and803(ip_12_35,x[12],y[35]);
and and804(ip_12_36,x[12],y[36]);
and and805(ip_12_37,x[12],y[37]);
and and806(ip_12_38,x[12],y[38]);
and and807(ip_12_39,x[12],y[39]);
and and808(ip_12_40,x[12],y[40]);
and and809(ip_12_41,x[12],y[41]);
and and810(ip_12_42,x[12],y[42]);
and and811(ip_12_43,x[12],y[43]);
and and812(ip_12_44,x[12],y[44]);
and and813(ip_12_45,x[12],y[45]);
and and814(ip_12_46,x[12],y[46]);
and and815(ip_12_47,x[12],y[47]);
and and816(ip_12_48,x[12],y[48]);
and and817(ip_12_49,x[12],y[49]);
and and818(ip_12_50,x[12],y[50]);
and and819(ip_12_51,x[12],y[51]);
and and820(ip_12_52,x[12],y[52]);
and and821(ip_12_53,x[12],y[53]);
and and822(ip_12_54,x[12],y[54]);
and and823(ip_12_55,x[12],y[55]);
and and824(ip_12_56,x[12],y[56]);
and and825(ip_12_57,x[12],y[57]);
and and826(ip_12_58,x[12],y[58]);
and and827(ip_12_59,x[12],y[59]);
and and828(ip_12_60,x[12],y[60]);
and and829(ip_12_61,x[12],y[61]);
and and830(ip_12_62,x[12],y[62]);
and and831(ip_12_63,x[12],y[63]);
and and832(ip_13_0,x[13],y[0]);
and and833(ip_13_1,x[13],y[1]);
and and834(ip_13_2,x[13],y[2]);
and and835(ip_13_3,x[13],y[3]);
and and836(ip_13_4,x[13],y[4]);
and and837(ip_13_5,x[13],y[5]);
and and838(ip_13_6,x[13],y[6]);
and and839(ip_13_7,x[13],y[7]);
and and840(ip_13_8,x[13],y[8]);
and and841(ip_13_9,x[13],y[9]);
and and842(ip_13_10,x[13],y[10]);
and and843(ip_13_11,x[13],y[11]);
and and844(ip_13_12,x[13],y[12]);
and and845(ip_13_13,x[13],y[13]);
and and846(ip_13_14,x[13],y[14]);
and and847(ip_13_15,x[13],y[15]);
and and848(ip_13_16,x[13],y[16]);
and and849(ip_13_17,x[13],y[17]);
and and850(ip_13_18,x[13],y[18]);
and and851(ip_13_19,x[13],y[19]);
and and852(ip_13_20,x[13],y[20]);
and and853(ip_13_21,x[13],y[21]);
and and854(ip_13_22,x[13],y[22]);
and and855(ip_13_23,x[13],y[23]);
and and856(ip_13_24,x[13],y[24]);
and and857(ip_13_25,x[13],y[25]);
and and858(ip_13_26,x[13],y[26]);
and and859(ip_13_27,x[13],y[27]);
and and860(ip_13_28,x[13],y[28]);
and and861(ip_13_29,x[13],y[29]);
and and862(ip_13_30,x[13],y[30]);
and and863(ip_13_31,x[13],y[31]);
and and864(ip_13_32,x[13],y[32]);
and and865(ip_13_33,x[13],y[33]);
and and866(ip_13_34,x[13],y[34]);
and and867(ip_13_35,x[13],y[35]);
and and868(ip_13_36,x[13],y[36]);
and and869(ip_13_37,x[13],y[37]);
and and870(ip_13_38,x[13],y[38]);
and and871(ip_13_39,x[13],y[39]);
and and872(ip_13_40,x[13],y[40]);
and and873(ip_13_41,x[13],y[41]);
and and874(ip_13_42,x[13],y[42]);
and and875(ip_13_43,x[13],y[43]);
and and876(ip_13_44,x[13],y[44]);
and and877(ip_13_45,x[13],y[45]);
and and878(ip_13_46,x[13],y[46]);
and and879(ip_13_47,x[13],y[47]);
and and880(ip_13_48,x[13],y[48]);
and and881(ip_13_49,x[13],y[49]);
and and882(ip_13_50,x[13],y[50]);
and and883(ip_13_51,x[13],y[51]);
and and884(ip_13_52,x[13],y[52]);
and and885(ip_13_53,x[13],y[53]);
and and886(ip_13_54,x[13],y[54]);
and and887(ip_13_55,x[13],y[55]);
and and888(ip_13_56,x[13],y[56]);
and and889(ip_13_57,x[13],y[57]);
and and890(ip_13_58,x[13],y[58]);
and and891(ip_13_59,x[13],y[59]);
and and892(ip_13_60,x[13],y[60]);
and and893(ip_13_61,x[13],y[61]);
and and894(ip_13_62,x[13],y[62]);
and and895(ip_13_63,x[13],y[63]);
and and896(ip_14_0,x[14],y[0]);
and and897(ip_14_1,x[14],y[1]);
and and898(ip_14_2,x[14],y[2]);
and and899(ip_14_3,x[14],y[3]);
and and900(ip_14_4,x[14],y[4]);
and and901(ip_14_5,x[14],y[5]);
and and902(ip_14_6,x[14],y[6]);
and and903(ip_14_7,x[14],y[7]);
and and904(ip_14_8,x[14],y[8]);
and and905(ip_14_9,x[14],y[9]);
and and906(ip_14_10,x[14],y[10]);
and and907(ip_14_11,x[14],y[11]);
and and908(ip_14_12,x[14],y[12]);
and and909(ip_14_13,x[14],y[13]);
and and910(ip_14_14,x[14],y[14]);
and and911(ip_14_15,x[14],y[15]);
and and912(ip_14_16,x[14],y[16]);
and and913(ip_14_17,x[14],y[17]);
and and914(ip_14_18,x[14],y[18]);
and and915(ip_14_19,x[14],y[19]);
and and916(ip_14_20,x[14],y[20]);
and and917(ip_14_21,x[14],y[21]);
and and918(ip_14_22,x[14],y[22]);
and and919(ip_14_23,x[14],y[23]);
and and920(ip_14_24,x[14],y[24]);
and and921(ip_14_25,x[14],y[25]);
and and922(ip_14_26,x[14],y[26]);
and and923(ip_14_27,x[14],y[27]);
and and924(ip_14_28,x[14],y[28]);
and and925(ip_14_29,x[14],y[29]);
and and926(ip_14_30,x[14],y[30]);
and and927(ip_14_31,x[14],y[31]);
and and928(ip_14_32,x[14],y[32]);
and and929(ip_14_33,x[14],y[33]);
and and930(ip_14_34,x[14],y[34]);
and and931(ip_14_35,x[14],y[35]);
and and932(ip_14_36,x[14],y[36]);
and and933(ip_14_37,x[14],y[37]);
and and934(ip_14_38,x[14],y[38]);
and and935(ip_14_39,x[14],y[39]);
and and936(ip_14_40,x[14],y[40]);
and and937(ip_14_41,x[14],y[41]);
and and938(ip_14_42,x[14],y[42]);
and and939(ip_14_43,x[14],y[43]);
and and940(ip_14_44,x[14],y[44]);
and and941(ip_14_45,x[14],y[45]);
and and942(ip_14_46,x[14],y[46]);
and and943(ip_14_47,x[14],y[47]);
and and944(ip_14_48,x[14],y[48]);
and and945(ip_14_49,x[14],y[49]);
and and946(ip_14_50,x[14],y[50]);
and and947(ip_14_51,x[14],y[51]);
and and948(ip_14_52,x[14],y[52]);
and and949(ip_14_53,x[14],y[53]);
and and950(ip_14_54,x[14],y[54]);
and and951(ip_14_55,x[14],y[55]);
and and952(ip_14_56,x[14],y[56]);
and and953(ip_14_57,x[14],y[57]);
and and954(ip_14_58,x[14],y[58]);
and and955(ip_14_59,x[14],y[59]);
and and956(ip_14_60,x[14],y[60]);
and and957(ip_14_61,x[14],y[61]);
and and958(ip_14_62,x[14],y[62]);
and and959(ip_14_63,x[14],y[63]);
and and960(ip_15_0,x[15],y[0]);
and and961(ip_15_1,x[15],y[1]);
and and962(ip_15_2,x[15],y[2]);
and and963(ip_15_3,x[15],y[3]);
and and964(ip_15_4,x[15],y[4]);
and and965(ip_15_5,x[15],y[5]);
and and966(ip_15_6,x[15],y[6]);
and and967(ip_15_7,x[15],y[7]);
and and968(ip_15_8,x[15],y[8]);
and and969(ip_15_9,x[15],y[9]);
and and970(ip_15_10,x[15],y[10]);
and and971(ip_15_11,x[15],y[11]);
and and972(ip_15_12,x[15],y[12]);
and and973(ip_15_13,x[15],y[13]);
and and974(ip_15_14,x[15],y[14]);
and and975(ip_15_15,x[15],y[15]);
and and976(ip_15_16,x[15],y[16]);
and and977(ip_15_17,x[15],y[17]);
and and978(ip_15_18,x[15],y[18]);
and and979(ip_15_19,x[15],y[19]);
and and980(ip_15_20,x[15],y[20]);
and and981(ip_15_21,x[15],y[21]);
and and982(ip_15_22,x[15],y[22]);
and and983(ip_15_23,x[15],y[23]);
and and984(ip_15_24,x[15],y[24]);
and and985(ip_15_25,x[15],y[25]);
and and986(ip_15_26,x[15],y[26]);
and and987(ip_15_27,x[15],y[27]);
and and988(ip_15_28,x[15],y[28]);
and and989(ip_15_29,x[15],y[29]);
and and990(ip_15_30,x[15],y[30]);
and and991(ip_15_31,x[15],y[31]);
and and992(ip_15_32,x[15],y[32]);
and and993(ip_15_33,x[15],y[33]);
and and994(ip_15_34,x[15],y[34]);
and and995(ip_15_35,x[15],y[35]);
and and996(ip_15_36,x[15],y[36]);
and and997(ip_15_37,x[15],y[37]);
and and998(ip_15_38,x[15],y[38]);
and and999(ip_15_39,x[15],y[39]);
and and1000(ip_15_40,x[15],y[40]);
and and1001(ip_15_41,x[15],y[41]);
and and1002(ip_15_42,x[15],y[42]);
and and1003(ip_15_43,x[15],y[43]);
and and1004(ip_15_44,x[15],y[44]);
and and1005(ip_15_45,x[15],y[45]);
and and1006(ip_15_46,x[15],y[46]);
and and1007(ip_15_47,x[15],y[47]);
and and1008(ip_15_48,x[15],y[48]);
and and1009(ip_15_49,x[15],y[49]);
and and1010(ip_15_50,x[15],y[50]);
and and1011(ip_15_51,x[15],y[51]);
and and1012(ip_15_52,x[15],y[52]);
and and1013(ip_15_53,x[15],y[53]);
and and1014(ip_15_54,x[15],y[54]);
and and1015(ip_15_55,x[15],y[55]);
and and1016(ip_15_56,x[15],y[56]);
and and1017(ip_15_57,x[15],y[57]);
and and1018(ip_15_58,x[15],y[58]);
and and1019(ip_15_59,x[15],y[59]);
and and1020(ip_15_60,x[15],y[60]);
and and1021(ip_15_61,x[15],y[61]);
and and1022(ip_15_62,x[15],y[62]);
and and1023(ip_15_63,x[15],y[63]);
and and1024(ip_16_0,x[16],y[0]);
and and1025(ip_16_1,x[16],y[1]);
and and1026(ip_16_2,x[16],y[2]);
and and1027(ip_16_3,x[16],y[3]);
and and1028(ip_16_4,x[16],y[4]);
and and1029(ip_16_5,x[16],y[5]);
and and1030(ip_16_6,x[16],y[6]);
and and1031(ip_16_7,x[16],y[7]);
and and1032(ip_16_8,x[16],y[8]);
and and1033(ip_16_9,x[16],y[9]);
and and1034(ip_16_10,x[16],y[10]);
and and1035(ip_16_11,x[16],y[11]);
and and1036(ip_16_12,x[16],y[12]);
and and1037(ip_16_13,x[16],y[13]);
and and1038(ip_16_14,x[16],y[14]);
and and1039(ip_16_15,x[16],y[15]);
and and1040(ip_16_16,x[16],y[16]);
and and1041(ip_16_17,x[16],y[17]);
and and1042(ip_16_18,x[16],y[18]);
and and1043(ip_16_19,x[16],y[19]);
and and1044(ip_16_20,x[16],y[20]);
and and1045(ip_16_21,x[16],y[21]);
and and1046(ip_16_22,x[16],y[22]);
and and1047(ip_16_23,x[16],y[23]);
and and1048(ip_16_24,x[16],y[24]);
and and1049(ip_16_25,x[16],y[25]);
and and1050(ip_16_26,x[16],y[26]);
and and1051(ip_16_27,x[16],y[27]);
and and1052(ip_16_28,x[16],y[28]);
and and1053(ip_16_29,x[16],y[29]);
and and1054(ip_16_30,x[16],y[30]);
and and1055(ip_16_31,x[16],y[31]);
and and1056(ip_16_32,x[16],y[32]);
and and1057(ip_16_33,x[16],y[33]);
and and1058(ip_16_34,x[16],y[34]);
and and1059(ip_16_35,x[16],y[35]);
and and1060(ip_16_36,x[16],y[36]);
and and1061(ip_16_37,x[16],y[37]);
and and1062(ip_16_38,x[16],y[38]);
and and1063(ip_16_39,x[16],y[39]);
and and1064(ip_16_40,x[16],y[40]);
and and1065(ip_16_41,x[16],y[41]);
and and1066(ip_16_42,x[16],y[42]);
and and1067(ip_16_43,x[16],y[43]);
and and1068(ip_16_44,x[16],y[44]);
and and1069(ip_16_45,x[16],y[45]);
and and1070(ip_16_46,x[16],y[46]);
and and1071(ip_16_47,x[16],y[47]);
and and1072(ip_16_48,x[16],y[48]);
and and1073(ip_16_49,x[16],y[49]);
and and1074(ip_16_50,x[16],y[50]);
and and1075(ip_16_51,x[16],y[51]);
and and1076(ip_16_52,x[16],y[52]);
and and1077(ip_16_53,x[16],y[53]);
and and1078(ip_16_54,x[16],y[54]);
and and1079(ip_16_55,x[16],y[55]);
and and1080(ip_16_56,x[16],y[56]);
and and1081(ip_16_57,x[16],y[57]);
and and1082(ip_16_58,x[16],y[58]);
and and1083(ip_16_59,x[16],y[59]);
and and1084(ip_16_60,x[16],y[60]);
and and1085(ip_16_61,x[16],y[61]);
and and1086(ip_16_62,x[16],y[62]);
and and1087(ip_16_63,x[16],y[63]);
and and1088(ip_17_0,x[17],y[0]);
and and1089(ip_17_1,x[17],y[1]);
and and1090(ip_17_2,x[17],y[2]);
and and1091(ip_17_3,x[17],y[3]);
and and1092(ip_17_4,x[17],y[4]);
and and1093(ip_17_5,x[17],y[5]);
and and1094(ip_17_6,x[17],y[6]);
and and1095(ip_17_7,x[17],y[7]);
and and1096(ip_17_8,x[17],y[8]);
and and1097(ip_17_9,x[17],y[9]);
and and1098(ip_17_10,x[17],y[10]);
and and1099(ip_17_11,x[17],y[11]);
and and1100(ip_17_12,x[17],y[12]);
and and1101(ip_17_13,x[17],y[13]);
and and1102(ip_17_14,x[17],y[14]);
and and1103(ip_17_15,x[17],y[15]);
and and1104(ip_17_16,x[17],y[16]);
and and1105(ip_17_17,x[17],y[17]);
and and1106(ip_17_18,x[17],y[18]);
and and1107(ip_17_19,x[17],y[19]);
and and1108(ip_17_20,x[17],y[20]);
and and1109(ip_17_21,x[17],y[21]);
and and1110(ip_17_22,x[17],y[22]);
and and1111(ip_17_23,x[17],y[23]);
and and1112(ip_17_24,x[17],y[24]);
and and1113(ip_17_25,x[17],y[25]);
and and1114(ip_17_26,x[17],y[26]);
and and1115(ip_17_27,x[17],y[27]);
and and1116(ip_17_28,x[17],y[28]);
and and1117(ip_17_29,x[17],y[29]);
and and1118(ip_17_30,x[17],y[30]);
and and1119(ip_17_31,x[17],y[31]);
and and1120(ip_17_32,x[17],y[32]);
and and1121(ip_17_33,x[17],y[33]);
and and1122(ip_17_34,x[17],y[34]);
and and1123(ip_17_35,x[17],y[35]);
and and1124(ip_17_36,x[17],y[36]);
and and1125(ip_17_37,x[17],y[37]);
and and1126(ip_17_38,x[17],y[38]);
and and1127(ip_17_39,x[17],y[39]);
and and1128(ip_17_40,x[17],y[40]);
and and1129(ip_17_41,x[17],y[41]);
and and1130(ip_17_42,x[17],y[42]);
and and1131(ip_17_43,x[17],y[43]);
and and1132(ip_17_44,x[17],y[44]);
and and1133(ip_17_45,x[17],y[45]);
and and1134(ip_17_46,x[17],y[46]);
and and1135(ip_17_47,x[17],y[47]);
and and1136(ip_17_48,x[17],y[48]);
and and1137(ip_17_49,x[17],y[49]);
and and1138(ip_17_50,x[17],y[50]);
and and1139(ip_17_51,x[17],y[51]);
and and1140(ip_17_52,x[17],y[52]);
and and1141(ip_17_53,x[17],y[53]);
and and1142(ip_17_54,x[17],y[54]);
and and1143(ip_17_55,x[17],y[55]);
and and1144(ip_17_56,x[17],y[56]);
and and1145(ip_17_57,x[17],y[57]);
and and1146(ip_17_58,x[17],y[58]);
and and1147(ip_17_59,x[17],y[59]);
and and1148(ip_17_60,x[17],y[60]);
and and1149(ip_17_61,x[17],y[61]);
and and1150(ip_17_62,x[17],y[62]);
and and1151(ip_17_63,x[17],y[63]);
and and1152(ip_18_0,x[18],y[0]);
and and1153(ip_18_1,x[18],y[1]);
and and1154(ip_18_2,x[18],y[2]);
and and1155(ip_18_3,x[18],y[3]);
and and1156(ip_18_4,x[18],y[4]);
and and1157(ip_18_5,x[18],y[5]);
and and1158(ip_18_6,x[18],y[6]);
and and1159(ip_18_7,x[18],y[7]);
and and1160(ip_18_8,x[18],y[8]);
and and1161(ip_18_9,x[18],y[9]);
and and1162(ip_18_10,x[18],y[10]);
and and1163(ip_18_11,x[18],y[11]);
and and1164(ip_18_12,x[18],y[12]);
and and1165(ip_18_13,x[18],y[13]);
and and1166(ip_18_14,x[18],y[14]);
and and1167(ip_18_15,x[18],y[15]);
and and1168(ip_18_16,x[18],y[16]);
and and1169(ip_18_17,x[18],y[17]);
and and1170(ip_18_18,x[18],y[18]);
and and1171(ip_18_19,x[18],y[19]);
and and1172(ip_18_20,x[18],y[20]);
and and1173(ip_18_21,x[18],y[21]);
and and1174(ip_18_22,x[18],y[22]);
and and1175(ip_18_23,x[18],y[23]);
and and1176(ip_18_24,x[18],y[24]);
and and1177(ip_18_25,x[18],y[25]);
and and1178(ip_18_26,x[18],y[26]);
and and1179(ip_18_27,x[18],y[27]);
and and1180(ip_18_28,x[18],y[28]);
and and1181(ip_18_29,x[18],y[29]);
and and1182(ip_18_30,x[18],y[30]);
and and1183(ip_18_31,x[18],y[31]);
and and1184(ip_18_32,x[18],y[32]);
and and1185(ip_18_33,x[18],y[33]);
and and1186(ip_18_34,x[18],y[34]);
and and1187(ip_18_35,x[18],y[35]);
and and1188(ip_18_36,x[18],y[36]);
and and1189(ip_18_37,x[18],y[37]);
and and1190(ip_18_38,x[18],y[38]);
and and1191(ip_18_39,x[18],y[39]);
and and1192(ip_18_40,x[18],y[40]);
and and1193(ip_18_41,x[18],y[41]);
and and1194(ip_18_42,x[18],y[42]);
and and1195(ip_18_43,x[18],y[43]);
and and1196(ip_18_44,x[18],y[44]);
and and1197(ip_18_45,x[18],y[45]);
and and1198(ip_18_46,x[18],y[46]);
and and1199(ip_18_47,x[18],y[47]);
and and1200(ip_18_48,x[18],y[48]);
and and1201(ip_18_49,x[18],y[49]);
and and1202(ip_18_50,x[18],y[50]);
and and1203(ip_18_51,x[18],y[51]);
and and1204(ip_18_52,x[18],y[52]);
and and1205(ip_18_53,x[18],y[53]);
and and1206(ip_18_54,x[18],y[54]);
and and1207(ip_18_55,x[18],y[55]);
and and1208(ip_18_56,x[18],y[56]);
and and1209(ip_18_57,x[18],y[57]);
and and1210(ip_18_58,x[18],y[58]);
and and1211(ip_18_59,x[18],y[59]);
and and1212(ip_18_60,x[18],y[60]);
and and1213(ip_18_61,x[18],y[61]);
and and1214(ip_18_62,x[18],y[62]);
and and1215(ip_18_63,x[18],y[63]);
and and1216(ip_19_0,x[19],y[0]);
and and1217(ip_19_1,x[19],y[1]);
and and1218(ip_19_2,x[19],y[2]);
and and1219(ip_19_3,x[19],y[3]);
and and1220(ip_19_4,x[19],y[4]);
and and1221(ip_19_5,x[19],y[5]);
and and1222(ip_19_6,x[19],y[6]);
and and1223(ip_19_7,x[19],y[7]);
and and1224(ip_19_8,x[19],y[8]);
and and1225(ip_19_9,x[19],y[9]);
and and1226(ip_19_10,x[19],y[10]);
and and1227(ip_19_11,x[19],y[11]);
and and1228(ip_19_12,x[19],y[12]);
and and1229(ip_19_13,x[19],y[13]);
and and1230(ip_19_14,x[19],y[14]);
and and1231(ip_19_15,x[19],y[15]);
and and1232(ip_19_16,x[19],y[16]);
and and1233(ip_19_17,x[19],y[17]);
and and1234(ip_19_18,x[19],y[18]);
and and1235(ip_19_19,x[19],y[19]);
and and1236(ip_19_20,x[19],y[20]);
and and1237(ip_19_21,x[19],y[21]);
and and1238(ip_19_22,x[19],y[22]);
and and1239(ip_19_23,x[19],y[23]);
and and1240(ip_19_24,x[19],y[24]);
and and1241(ip_19_25,x[19],y[25]);
and and1242(ip_19_26,x[19],y[26]);
and and1243(ip_19_27,x[19],y[27]);
and and1244(ip_19_28,x[19],y[28]);
and and1245(ip_19_29,x[19],y[29]);
and and1246(ip_19_30,x[19],y[30]);
and and1247(ip_19_31,x[19],y[31]);
and and1248(ip_19_32,x[19],y[32]);
and and1249(ip_19_33,x[19],y[33]);
and and1250(ip_19_34,x[19],y[34]);
and and1251(ip_19_35,x[19],y[35]);
and and1252(ip_19_36,x[19],y[36]);
and and1253(ip_19_37,x[19],y[37]);
and and1254(ip_19_38,x[19],y[38]);
and and1255(ip_19_39,x[19],y[39]);
and and1256(ip_19_40,x[19],y[40]);
and and1257(ip_19_41,x[19],y[41]);
and and1258(ip_19_42,x[19],y[42]);
and and1259(ip_19_43,x[19],y[43]);
and and1260(ip_19_44,x[19],y[44]);
and and1261(ip_19_45,x[19],y[45]);
and and1262(ip_19_46,x[19],y[46]);
and and1263(ip_19_47,x[19],y[47]);
and and1264(ip_19_48,x[19],y[48]);
and and1265(ip_19_49,x[19],y[49]);
and and1266(ip_19_50,x[19],y[50]);
and and1267(ip_19_51,x[19],y[51]);
and and1268(ip_19_52,x[19],y[52]);
and and1269(ip_19_53,x[19],y[53]);
and and1270(ip_19_54,x[19],y[54]);
and and1271(ip_19_55,x[19],y[55]);
and and1272(ip_19_56,x[19],y[56]);
and and1273(ip_19_57,x[19],y[57]);
and and1274(ip_19_58,x[19],y[58]);
and and1275(ip_19_59,x[19],y[59]);
and and1276(ip_19_60,x[19],y[60]);
and and1277(ip_19_61,x[19],y[61]);
and and1278(ip_19_62,x[19],y[62]);
and and1279(ip_19_63,x[19],y[63]);
and and1280(ip_20_0,x[20],y[0]);
and and1281(ip_20_1,x[20],y[1]);
and and1282(ip_20_2,x[20],y[2]);
and and1283(ip_20_3,x[20],y[3]);
and and1284(ip_20_4,x[20],y[4]);
and and1285(ip_20_5,x[20],y[5]);
and and1286(ip_20_6,x[20],y[6]);
and and1287(ip_20_7,x[20],y[7]);
and and1288(ip_20_8,x[20],y[8]);
and and1289(ip_20_9,x[20],y[9]);
and and1290(ip_20_10,x[20],y[10]);
and and1291(ip_20_11,x[20],y[11]);
and and1292(ip_20_12,x[20],y[12]);
and and1293(ip_20_13,x[20],y[13]);
and and1294(ip_20_14,x[20],y[14]);
and and1295(ip_20_15,x[20],y[15]);
and and1296(ip_20_16,x[20],y[16]);
and and1297(ip_20_17,x[20],y[17]);
and and1298(ip_20_18,x[20],y[18]);
and and1299(ip_20_19,x[20],y[19]);
and and1300(ip_20_20,x[20],y[20]);
and and1301(ip_20_21,x[20],y[21]);
and and1302(ip_20_22,x[20],y[22]);
and and1303(ip_20_23,x[20],y[23]);
and and1304(ip_20_24,x[20],y[24]);
and and1305(ip_20_25,x[20],y[25]);
and and1306(ip_20_26,x[20],y[26]);
and and1307(ip_20_27,x[20],y[27]);
and and1308(ip_20_28,x[20],y[28]);
and and1309(ip_20_29,x[20],y[29]);
and and1310(ip_20_30,x[20],y[30]);
and and1311(ip_20_31,x[20],y[31]);
and and1312(ip_20_32,x[20],y[32]);
and and1313(ip_20_33,x[20],y[33]);
and and1314(ip_20_34,x[20],y[34]);
and and1315(ip_20_35,x[20],y[35]);
and and1316(ip_20_36,x[20],y[36]);
and and1317(ip_20_37,x[20],y[37]);
and and1318(ip_20_38,x[20],y[38]);
and and1319(ip_20_39,x[20],y[39]);
and and1320(ip_20_40,x[20],y[40]);
and and1321(ip_20_41,x[20],y[41]);
and and1322(ip_20_42,x[20],y[42]);
and and1323(ip_20_43,x[20],y[43]);
and and1324(ip_20_44,x[20],y[44]);
and and1325(ip_20_45,x[20],y[45]);
and and1326(ip_20_46,x[20],y[46]);
and and1327(ip_20_47,x[20],y[47]);
and and1328(ip_20_48,x[20],y[48]);
and and1329(ip_20_49,x[20],y[49]);
and and1330(ip_20_50,x[20],y[50]);
and and1331(ip_20_51,x[20],y[51]);
and and1332(ip_20_52,x[20],y[52]);
and and1333(ip_20_53,x[20],y[53]);
and and1334(ip_20_54,x[20],y[54]);
and and1335(ip_20_55,x[20],y[55]);
and and1336(ip_20_56,x[20],y[56]);
and and1337(ip_20_57,x[20],y[57]);
and and1338(ip_20_58,x[20],y[58]);
and and1339(ip_20_59,x[20],y[59]);
and and1340(ip_20_60,x[20],y[60]);
and and1341(ip_20_61,x[20],y[61]);
and and1342(ip_20_62,x[20],y[62]);
and and1343(ip_20_63,x[20],y[63]);
and and1344(ip_21_0,x[21],y[0]);
and and1345(ip_21_1,x[21],y[1]);
and and1346(ip_21_2,x[21],y[2]);
and and1347(ip_21_3,x[21],y[3]);
and and1348(ip_21_4,x[21],y[4]);
and and1349(ip_21_5,x[21],y[5]);
and and1350(ip_21_6,x[21],y[6]);
and and1351(ip_21_7,x[21],y[7]);
and and1352(ip_21_8,x[21],y[8]);
and and1353(ip_21_9,x[21],y[9]);
and and1354(ip_21_10,x[21],y[10]);
and and1355(ip_21_11,x[21],y[11]);
and and1356(ip_21_12,x[21],y[12]);
and and1357(ip_21_13,x[21],y[13]);
and and1358(ip_21_14,x[21],y[14]);
and and1359(ip_21_15,x[21],y[15]);
and and1360(ip_21_16,x[21],y[16]);
and and1361(ip_21_17,x[21],y[17]);
and and1362(ip_21_18,x[21],y[18]);
and and1363(ip_21_19,x[21],y[19]);
and and1364(ip_21_20,x[21],y[20]);
and and1365(ip_21_21,x[21],y[21]);
and and1366(ip_21_22,x[21],y[22]);
and and1367(ip_21_23,x[21],y[23]);
and and1368(ip_21_24,x[21],y[24]);
and and1369(ip_21_25,x[21],y[25]);
and and1370(ip_21_26,x[21],y[26]);
and and1371(ip_21_27,x[21],y[27]);
and and1372(ip_21_28,x[21],y[28]);
and and1373(ip_21_29,x[21],y[29]);
and and1374(ip_21_30,x[21],y[30]);
and and1375(ip_21_31,x[21],y[31]);
and and1376(ip_21_32,x[21],y[32]);
and and1377(ip_21_33,x[21],y[33]);
and and1378(ip_21_34,x[21],y[34]);
and and1379(ip_21_35,x[21],y[35]);
and and1380(ip_21_36,x[21],y[36]);
and and1381(ip_21_37,x[21],y[37]);
and and1382(ip_21_38,x[21],y[38]);
and and1383(ip_21_39,x[21],y[39]);
and and1384(ip_21_40,x[21],y[40]);
and and1385(ip_21_41,x[21],y[41]);
and and1386(ip_21_42,x[21],y[42]);
and and1387(ip_21_43,x[21],y[43]);
and and1388(ip_21_44,x[21],y[44]);
and and1389(ip_21_45,x[21],y[45]);
and and1390(ip_21_46,x[21],y[46]);
and and1391(ip_21_47,x[21],y[47]);
and and1392(ip_21_48,x[21],y[48]);
and and1393(ip_21_49,x[21],y[49]);
and and1394(ip_21_50,x[21],y[50]);
and and1395(ip_21_51,x[21],y[51]);
and and1396(ip_21_52,x[21],y[52]);
and and1397(ip_21_53,x[21],y[53]);
and and1398(ip_21_54,x[21],y[54]);
and and1399(ip_21_55,x[21],y[55]);
and and1400(ip_21_56,x[21],y[56]);
and and1401(ip_21_57,x[21],y[57]);
and and1402(ip_21_58,x[21],y[58]);
and and1403(ip_21_59,x[21],y[59]);
and and1404(ip_21_60,x[21],y[60]);
and and1405(ip_21_61,x[21],y[61]);
and and1406(ip_21_62,x[21],y[62]);
and and1407(ip_21_63,x[21],y[63]);
and and1408(ip_22_0,x[22],y[0]);
and and1409(ip_22_1,x[22],y[1]);
and and1410(ip_22_2,x[22],y[2]);
and and1411(ip_22_3,x[22],y[3]);
and and1412(ip_22_4,x[22],y[4]);
and and1413(ip_22_5,x[22],y[5]);
and and1414(ip_22_6,x[22],y[6]);
and and1415(ip_22_7,x[22],y[7]);
and and1416(ip_22_8,x[22],y[8]);
and and1417(ip_22_9,x[22],y[9]);
and and1418(ip_22_10,x[22],y[10]);
and and1419(ip_22_11,x[22],y[11]);
and and1420(ip_22_12,x[22],y[12]);
and and1421(ip_22_13,x[22],y[13]);
and and1422(ip_22_14,x[22],y[14]);
and and1423(ip_22_15,x[22],y[15]);
and and1424(ip_22_16,x[22],y[16]);
and and1425(ip_22_17,x[22],y[17]);
and and1426(ip_22_18,x[22],y[18]);
and and1427(ip_22_19,x[22],y[19]);
and and1428(ip_22_20,x[22],y[20]);
and and1429(ip_22_21,x[22],y[21]);
and and1430(ip_22_22,x[22],y[22]);
and and1431(ip_22_23,x[22],y[23]);
and and1432(ip_22_24,x[22],y[24]);
and and1433(ip_22_25,x[22],y[25]);
and and1434(ip_22_26,x[22],y[26]);
and and1435(ip_22_27,x[22],y[27]);
and and1436(ip_22_28,x[22],y[28]);
and and1437(ip_22_29,x[22],y[29]);
and and1438(ip_22_30,x[22],y[30]);
and and1439(ip_22_31,x[22],y[31]);
and and1440(ip_22_32,x[22],y[32]);
and and1441(ip_22_33,x[22],y[33]);
and and1442(ip_22_34,x[22],y[34]);
and and1443(ip_22_35,x[22],y[35]);
and and1444(ip_22_36,x[22],y[36]);
and and1445(ip_22_37,x[22],y[37]);
and and1446(ip_22_38,x[22],y[38]);
and and1447(ip_22_39,x[22],y[39]);
and and1448(ip_22_40,x[22],y[40]);
and and1449(ip_22_41,x[22],y[41]);
and and1450(ip_22_42,x[22],y[42]);
and and1451(ip_22_43,x[22],y[43]);
and and1452(ip_22_44,x[22],y[44]);
and and1453(ip_22_45,x[22],y[45]);
and and1454(ip_22_46,x[22],y[46]);
and and1455(ip_22_47,x[22],y[47]);
and and1456(ip_22_48,x[22],y[48]);
and and1457(ip_22_49,x[22],y[49]);
and and1458(ip_22_50,x[22],y[50]);
and and1459(ip_22_51,x[22],y[51]);
and and1460(ip_22_52,x[22],y[52]);
and and1461(ip_22_53,x[22],y[53]);
and and1462(ip_22_54,x[22],y[54]);
and and1463(ip_22_55,x[22],y[55]);
and and1464(ip_22_56,x[22],y[56]);
and and1465(ip_22_57,x[22],y[57]);
and and1466(ip_22_58,x[22],y[58]);
and and1467(ip_22_59,x[22],y[59]);
and and1468(ip_22_60,x[22],y[60]);
and and1469(ip_22_61,x[22],y[61]);
and and1470(ip_22_62,x[22],y[62]);
and and1471(ip_22_63,x[22],y[63]);
and and1472(ip_23_0,x[23],y[0]);
and and1473(ip_23_1,x[23],y[1]);
and and1474(ip_23_2,x[23],y[2]);
and and1475(ip_23_3,x[23],y[3]);
and and1476(ip_23_4,x[23],y[4]);
and and1477(ip_23_5,x[23],y[5]);
and and1478(ip_23_6,x[23],y[6]);
and and1479(ip_23_7,x[23],y[7]);
and and1480(ip_23_8,x[23],y[8]);
and and1481(ip_23_9,x[23],y[9]);
and and1482(ip_23_10,x[23],y[10]);
and and1483(ip_23_11,x[23],y[11]);
and and1484(ip_23_12,x[23],y[12]);
and and1485(ip_23_13,x[23],y[13]);
and and1486(ip_23_14,x[23],y[14]);
and and1487(ip_23_15,x[23],y[15]);
and and1488(ip_23_16,x[23],y[16]);
and and1489(ip_23_17,x[23],y[17]);
and and1490(ip_23_18,x[23],y[18]);
and and1491(ip_23_19,x[23],y[19]);
and and1492(ip_23_20,x[23],y[20]);
and and1493(ip_23_21,x[23],y[21]);
and and1494(ip_23_22,x[23],y[22]);
and and1495(ip_23_23,x[23],y[23]);
and and1496(ip_23_24,x[23],y[24]);
and and1497(ip_23_25,x[23],y[25]);
and and1498(ip_23_26,x[23],y[26]);
and and1499(ip_23_27,x[23],y[27]);
and and1500(ip_23_28,x[23],y[28]);
and and1501(ip_23_29,x[23],y[29]);
and and1502(ip_23_30,x[23],y[30]);
and and1503(ip_23_31,x[23],y[31]);
and and1504(ip_23_32,x[23],y[32]);
and and1505(ip_23_33,x[23],y[33]);
and and1506(ip_23_34,x[23],y[34]);
and and1507(ip_23_35,x[23],y[35]);
and and1508(ip_23_36,x[23],y[36]);
and and1509(ip_23_37,x[23],y[37]);
and and1510(ip_23_38,x[23],y[38]);
and and1511(ip_23_39,x[23],y[39]);
and and1512(ip_23_40,x[23],y[40]);
and and1513(ip_23_41,x[23],y[41]);
and and1514(ip_23_42,x[23],y[42]);
and and1515(ip_23_43,x[23],y[43]);
and and1516(ip_23_44,x[23],y[44]);
and and1517(ip_23_45,x[23],y[45]);
and and1518(ip_23_46,x[23],y[46]);
and and1519(ip_23_47,x[23],y[47]);
and and1520(ip_23_48,x[23],y[48]);
and and1521(ip_23_49,x[23],y[49]);
and and1522(ip_23_50,x[23],y[50]);
and and1523(ip_23_51,x[23],y[51]);
and and1524(ip_23_52,x[23],y[52]);
and and1525(ip_23_53,x[23],y[53]);
and and1526(ip_23_54,x[23],y[54]);
and and1527(ip_23_55,x[23],y[55]);
and and1528(ip_23_56,x[23],y[56]);
and and1529(ip_23_57,x[23],y[57]);
and and1530(ip_23_58,x[23],y[58]);
and and1531(ip_23_59,x[23],y[59]);
and and1532(ip_23_60,x[23],y[60]);
and and1533(ip_23_61,x[23],y[61]);
and and1534(ip_23_62,x[23],y[62]);
and and1535(ip_23_63,x[23],y[63]);
and and1536(ip_24_0,x[24],y[0]);
and and1537(ip_24_1,x[24],y[1]);
and and1538(ip_24_2,x[24],y[2]);
and and1539(ip_24_3,x[24],y[3]);
and and1540(ip_24_4,x[24],y[4]);
and and1541(ip_24_5,x[24],y[5]);
and and1542(ip_24_6,x[24],y[6]);
and and1543(ip_24_7,x[24],y[7]);
and and1544(ip_24_8,x[24],y[8]);
and and1545(ip_24_9,x[24],y[9]);
and and1546(ip_24_10,x[24],y[10]);
and and1547(ip_24_11,x[24],y[11]);
and and1548(ip_24_12,x[24],y[12]);
and and1549(ip_24_13,x[24],y[13]);
and and1550(ip_24_14,x[24],y[14]);
and and1551(ip_24_15,x[24],y[15]);
and and1552(ip_24_16,x[24],y[16]);
and and1553(ip_24_17,x[24],y[17]);
and and1554(ip_24_18,x[24],y[18]);
and and1555(ip_24_19,x[24],y[19]);
and and1556(ip_24_20,x[24],y[20]);
and and1557(ip_24_21,x[24],y[21]);
and and1558(ip_24_22,x[24],y[22]);
and and1559(ip_24_23,x[24],y[23]);
and and1560(ip_24_24,x[24],y[24]);
and and1561(ip_24_25,x[24],y[25]);
and and1562(ip_24_26,x[24],y[26]);
and and1563(ip_24_27,x[24],y[27]);
and and1564(ip_24_28,x[24],y[28]);
and and1565(ip_24_29,x[24],y[29]);
and and1566(ip_24_30,x[24],y[30]);
and and1567(ip_24_31,x[24],y[31]);
and and1568(ip_24_32,x[24],y[32]);
and and1569(ip_24_33,x[24],y[33]);
and and1570(ip_24_34,x[24],y[34]);
and and1571(ip_24_35,x[24],y[35]);
and and1572(ip_24_36,x[24],y[36]);
and and1573(ip_24_37,x[24],y[37]);
and and1574(ip_24_38,x[24],y[38]);
and and1575(ip_24_39,x[24],y[39]);
and and1576(ip_24_40,x[24],y[40]);
and and1577(ip_24_41,x[24],y[41]);
and and1578(ip_24_42,x[24],y[42]);
and and1579(ip_24_43,x[24],y[43]);
and and1580(ip_24_44,x[24],y[44]);
and and1581(ip_24_45,x[24],y[45]);
and and1582(ip_24_46,x[24],y[46]);
and and1583(ip_24_47,x[24],y[47]);
and and1584(ip_24_48,x[24],y[48]);
and and1585(ip_24_49,x[24],y[49]);
and and1586(ip_24_50,x[24],y[50]);
and and1587(ip_24_51,x[24],y[51]);
and and1588(ip_24_52,x[24],y[52]);
and and1589(ip_24_53,x[24],y[53]);
and and1590(ip_24_54,x[24],y[54]);
and and1591(ip_24_55,x[24],y[55]);
and and1592(ip_24_56,x[24],y[56]);
and and1593(ip_24_57,x[24],y[57]);
and and1594(ip_24_58,x[24],y[58]);
and and1595(ip_24_59,x[24],y[59]);
and and1596(ip_24_60,x[24],y[60]);
and and1597(ip_24_61,x[24],y[61]);
and and1598(ip_24_62,x[24],y[62]);
and and1599(ip_24_63,x[24],y[63]);
and and1600(ip_25_0,x[25],y[0]);
and and1601(ip_25_1,x[25],y[1]);
and and1602(ip_25_2,x[25],y[2]);
and and1603(ip_25_3,x[25],y[3]);
and and1604(ip_25_4,x[25],y[4]);
and and1605(ip_25_5,x[25],y[5]);
and and1606(ip_25_6,x[25],y[6]);
and and1607(ip_25_7,x[25],y[7]);
and and1608(ip_25_8,x[25],y[8]);
and and1609(ip_25_9,x[25],y[9]);
and and1610(ip_25_10,x[25],y[10]);
and and1611(ip_25_11,x[25],y[11]);
and and1612(ip_25_12,x[25],y[12]);
and and1613(ip_25_13,x[25],y[13]);
and and1614(ip_25_14,x[25],y[14]);
and and1615(ip_25_15,x[25],y[15]);
and and1616(ip_25_16,x[25],y[16]);
and and1617(ip_25_17,x[25],y[17]);
and and1618(ip_25_18,x[25],y[18]);
and and1619(ip_25_19,x[25],y[19]);
and and1620(ip_25_20,x[25],y[20]);
and and1621(ip_25_21,x[25],y[21]);
and and1622(ip_25_22,x[25],y[22]);
and and1623(ip_25_23,x[25],y[23]);
and and1624(ip_25_24,x[25],y[24]);
and and1625(ip_25_25,x[25],y[25]);
and and1626(ip_25_26,x[25],y[26]);
and and1627(ip_25_27,x[25],y[27]);
and and1628(ip_25_28,x[25],y[28]);
and and1629(ip_25_29,x[25],y[29]);
and and1630(ip_25_30,x[25],y[30]);
and and1631(ip_25_31,x[25],y[31]);
and and1632(ip_25_32,x[25],y[32]);
and and1633(ip_25_33,x[25],y[33]);
and and1634(ip_25_34,x[25],y[34]);
and and1635(ip_25_35,x[25],y[35]);
and and1636(ip_25_36,x[25],y[36]);
and and1637(ip_25_37,x[25],y[37]);
and and1638(ip_25_38,x[25],y[38]);
and and1639(ip_25_39,x[25],y[39]);
and and1640(ip_25_40,x[25],y[40]);
and and1641(ip_25_41,x[25],y[41]);
and and1642(ip_25_42,x[25],y[42]);
and and1643(ip_25_43,x[25],y[43]);
and and1644(ip_25_44,x[25],y[44]);
and and1645(ip_25_45,x[25],y[45]);
and and1646(ip_25_46,x[25],y[46]);
and and1647(ip_25_47,x[25],y[47]);
and and1648(ip_25_48,x[25],y[48]);
and and1649(ip_25_49,x[25],y[49]);
and and1650(ip_25_50,x[25],y[50]);
and and1651(ip_25_51,x[25],y[51]);
and and1652(ip_25_52,x[25],y[52]);
and and1653(ip_25_53,x[25],y[53]);
and and1654(ip_25_54,x[25],y[54]);
and and1655(ip_25_55,x[25],y[55]);
and and1656(ip_25_56,x[25],y[56]);
and and1657(ip_25_57,x[25],y[57]);
and and1658(ip_25_58,x[25],y[58]);
and and1659(ip_25_59,x[25],y[59]);
and and1660(ip_25_60,x[25],y[60]);
and and1661(ip_25_61,x[25],y[61]);
and and1662(ip_25_62,x[25],y[62]);
and and1663(ip_25_63,x[25],y[63]);
and and1664(ip_26_0,x[26],y[0]);
and and1665(ip_26_1,x[26],y[1]);
and and1666(ip_26_2,x[26],y[2]);
and and1667(ip_26_3,x[26],y[3]);
and and1668(ip_26_4,x[26],y[4]);
and and1669(ip_26_5,x[26],y[5]);
and and1670(ip_26_6,x[26],y[6]);
and and1671(ip_26_7,x[26],y[7]);
and and1672(ip_26_8,x[26],y[8]);
and and1673(ip_26_9,x[26],y[9]);
and and1674(ip_26_10,x[26],y[10]);
and and1675(ip_26_11,x[26],y[11]);
and and1676(ip_26_12,x[26],y[12]);
and and1677(ip_26_13,x[26],y[13]);
and and1678(ip_26_14,x[26],y[14]);
and and1679(ip_26_15,x[26],y[15]);
and and1680(ip_26_16,x[26],y[16]);
and and1681(ip_26_17,x[26],y[17]);
and and1682(ip_26_18,x[26],y[18]);
and and1683(ip_26_19,x[26],y[19]);
and and1684(ip_26_20,x[26],y[20]);
and and1685(ip_26_21,x[26],y[21]);
and and1686(ip_26_22,x[26],y[22]);
and and1687(ip_26_23,x[26],y[23]);
and and1688(ip_26_24,x[26],y[24]);
and and1689(ip_26_25,x[26],y[25]);
and and1690(ip_26_26,x[26],y[26]);
and and1691(ip_26_27,x[26],y[27]);
and and1692(ip_26_28,x[26],y[28]);
and and1693(ip_26_29,x[26],y[29]);
and and1694(ip_26_30,x[26],y[30]);
and and1695(ip_26_31,x[26],y[31]);
and and1696(ip_26_32,x[26],y[32]);
and and1697(ip_26_33,x[26],y[33]);
and and1698(ip_26_34,x[26],y[34]);
and and1699(ip_26_35,x[26],y[35]);
and and1700(ip_26_36,x[26],y[36]);
and and1701(ip_26_37,x[26],y[37]);
and and1702(ip_26_38,x[26],y[38]);
and and1703(ip_26_39,x[26],y[39]);
and and1704(ip_26_40,x[26],y[40]);
and and1705(ip_26_41,x[26],y[41]);
and and1706(ip_26_42,x[26],y[42]);
and and1707(ip_26_43,x[26],y[43]);
and and1708(ip_26_44,x[26],y[44]);
and and1709(ip_26_45,x[26],y[45]);
and and1710(ip_26_46,x[26],y[46]);
and and1711(ip_26_47,x[26],y[47]);
and and1712(ip_26_48,x[26],y[48]);
and and1713(ip_26_49,x[26],y[49]);
and and1714(ip_26_50,x[26],y[50]);
and and1715(ip_26_51,x[26],y[51]);
and and1716(ip_26_52,x[26],y[52]);
and and1717(ip_26_53,x[26],y[53]);
and and1718(ip_26_54,x[26],y[54]);
and and1719(ip_26_55,x[26],y[55]);
and and1720(ip_26_56,x[26],y[56]);
and and1721(ip_26_57,x[26],y[57]);
and and1722(ip_26_58,x[26],y[58]);
and and1723(ip_26_59,x[26],y[59]);
and and1724(ip_26_60,x[26],y[60]);
and and1725(ip_26_61,x[26],y[61]);
and and1726(ip_26_62,x[26],y[62]);
and and1727(ip_26_63,x[26],y[63]);
and and1728(ip_27_0,x[27],y[0]);
and and1729(ip_27_1,x[27],y[1]);
and and1730(ip_27_2,x[27],y[2]);
and and1731(ip_27_3,x[27],y[3]);
and and1732(ip_27_4,x[27],y[4]);
and and1733(ip_27_5,x[27],y[5]);
and and1734(ip_27_6,x[27],y[6]);
and and1735(ip_27_7,x[27],y[7]);
and and1736(ip_27_8,x[27],y[8]);
and and1737(ip_27_9,x[27],y[9]);
and and1738(ip_27_10,x[27],y[10]);
and and1739(ip_27_11,x[27],y[11]);
and and1740(ip_27_12,x[27],y[12]);
and and1741(ip_27_13,x[27],y[13]);
and and1742(ip_27_14,x[27],y[14]);
and and1743(ip_27_15,x[27],y[15]);
and and1744(ip_27_16,x[27],y[16]);
and and1745(ip_27_17,x[27],y[17]);
and and1746(ip_27_18,x[27],y[18]);
and and1747(ip_27_19,x[27],y[19]);
and and1748(ip_27_20,x[27],y[20]);
and and1749(ip_27_21,x[27],y[21]);
and and1750(ip_27_22,x[27],y[22]);
and and1751(ip_27_23,x[27],y[23]);
and and1752(ip_27_24,x[27],y[24]);
and and1753(ip_27_25,x[27],y[25]);
and and1754(ip_27_26,x[27],y[26]);
and and1755(ip_27_27,x[27],y[27]);
and and1756(ip_27_28,x[27],y[28]);
and and1757(ip_27_29,x[27],y[29]);
and and1758(ip_27_30,x[27],y[30]);
and and1759(ip_27_31,x[27],y[31]);
and and1760(ip_27_32,x[27],y[32]);
and and1761(ip_27_33,x[27],y[33]);
and and1762(ip_27_34,x[27],y[34]);
and and1763(ip_27_35,x[27],y[35]);
and and1764(ip_27_36,x[27],y[36]);
and and1765(ip_27_37,x[27],y[37]);
and and1766(ip_27_38,x[27],y[38]);
and and1767(ip_27_39,x[27],y[39]);
and and1768(ip_27_40,x[27],y[40]);
and and1769(ip_27_41,x[27],y[41]);
and and1770(ip_27_42,x[27],y[42]);
and and1771(ip_27_43,x[27],y[43]);
and and1772(ip_27_44,x[27],y[44]);
and and1773(ip_27_45,x[27],y[45]);
and and1774(ip_27_46,x[27],y[46]);
and and1775(ip_27_47,x[27],y[47]);
and and1776(ip_27_48,x[27],y[48]);
and and1777(ip_27_49,x[27],y[49]);
and and1778(ip_27_50,x[27],y[50]);
and and1779(ip_27_51,x[27],y[51]);
and and1780(ip_27_52,x[27],y[52]);
and and1781(ip_27_53,x[27],y[53]);
and and1782(ip_27_54,x[27],y[54]);
and and1783(ip_27_55,x[27],y[55]);
and and1784(ip_27_56,x[27],y[56]);
and and1785(ip_27_57,x[27],y[57]);
and and1786(ip_27_58,x[27],y[58]);
and and1787(ip_27_59,x[27],y[59]);
and and1788(ip_27_60,x[27],y[60]);
and and1789(ip_27_61,x[27],y[61]);
and and1790(ip_27_62,x[27],y[62]);
and and1791(ip_27_63,x[27],y[63]);
and and1792(ip_28_0,x[28],y[0]);
and and1793(ip_28_1,x[28],y[1]);
and and1794(ip_28_2,x[28],y[2]);
and and1795(ip_28_3,x[28],y[3]);
and and1796(ip_28_4,x[28],y[4]);
and and1797(ip_28_5,x[28],y[5]);
and and1798(ip_28_6,x[28],y[6]);
and and1799(ip_28_7,x[28],y[7]);
and and1800(ip_28_8,x[28],y[8]);
and and1801(ip_28_9,x[28],y[9]);
and and1802(ip_28_10,x[28],y[10]);
and and1803(ip_28_11,x[28],y[11]);
and and1804(ip_28_12,x[28],y[12]);
and and1805(ip_28_13,x[28],y[13]);
and and1806(ip_28_14,x[28],y[14]);
and and1807(ip_28_15,x[28],y[15]);
and and1808(ip_28_16,x[28],y[16]);
and and1809(ip_28_17,x[28],y[17]);
and and1810(ip_28_18,x[28],y[18]);
and and1811(ip_28_19,x[28],y[19]);
and and1812(ip_28_20,x[28],y[20]);
and and1813(ip_28_21,x[28],y[21]);
and and1814(ip_28_22,x[28],y[22]);
and and1815(ip_28_23,x[28],y[23]);
and and1816(ip_28_24,x[28],y[24]);
and and1817(ip_28_25,x[28],y[25]);
and and1818(ip_28_26,x[28],y[26]);
and and1819(ip_28_27,x[28],y[27]);
and and1820(ip_28_28,x[28],y[28]);
and and1821(ip_28_29,x[28],y[29]);
and and1822(ip_28_30,x[28],y[30]);
and and1823(ip_28_31,x[28],y[31]);
and and1824(ip_28_32,x[28],y[32]);
and and1825(ip_28_33,x[28],y[33]);
and and1826(ip_28_34,x[28],y[34]);
and and1827(ip_28_35,x[28],y[35]);
and and1828(ip_28_36,x[28],y[36]);
and and1829(ip_28_37,x[28],y[37]);
and and1830(ip_28_38,x[28],y[38]);
and and1831(ip_28_39,x[28],y[39]);
and and1832(ip_28_40,x[28],y[40]);
and and1833(ip_28_41,x[28],y[41]);
and and1834(ip_28_42,x[28],y[42]);
and and1835(ip_28_43,x[28],y[43]);
and and1836(ip_28_44,x[28],y[44]);
and and1837(ip_28_45,x[28],y[45]);
and and1838(ip_28_46,x[28],y[46]);
and and1839(ip_28_47,x[28],y[47]);
and and1840(ip_28_48,x[28],y[48]);
and and1841(ip_28_49,x[28],y[49]);
and and1842(ip_28_50,x[28],y[50]);
and and1843(ip_28_51,x[28],y[51]);
and and1844(ip_28_52,x[28],y[52]);
and and1845(ip_28_53,x[28],y[53]);
and and1846(ip_28_54,x[28],y[54]);
and and1847(ip_28_55,x[28],y[55]);
and and1848(ip_28_56,x[28],y[56]);
and and1849(ip_28_57,x[28],y[57]);
and and1850(ip_28_58,x[28],y[58]);
and and1851(ip_28_59,x[28],y[59]);
and and1852(ip_28_60,x[28],y[60]);
and and1853(ip_28_61,x[28],y[61]);
and and1854(ip_28_62,x[28],y[62]);
and and1855(ip_28_63,x[28],y[63]);
and and1856(ip_29_0,x[29],y[0]);
and and1857(ip_29_1,x[29],y[1]);
and and1858(ip_29_2,x[29],y[2]);
and and1859(ip_29_3,x[29],y[3]);
and and1860(ip_29_4,x[29],y[4]);
and and1861(ip_29_5,x[29],y[5]);
and and1862(ip_29_6,x[29],y[6]);
and and1863(ip_29_7,x[29],y[7]);
and and1864(ip_29_8,x[29],y[8]);
and and1865(ip_29_9,x[29],y[9]);
and and1866(ip_29_10,x[29],y[10]);
and and1867(ip_29_11,x[29],y[11]);
and and1868(ip_29_12,x[29],y[12]);
and and1869(ip_29_13,x[29],y[13]);
and and1870(ip_29_14,x[29],y[14]);
and and1871(ip_29_15,x[29],y[15]);
and and1872(ip_29_16,x[29],y[16]);
and and1873(ip_29_17,x[29],y[17]);
and and1874(ip_29_18,x[29],y[18]);
and and1875(ip_29_19,x[29],y[19]);
and and1876(ip_29_20,x[29],y[20]);
and and1877(ip_29_21,x[29],y[21]);
and and1878(ip_29_22,x[29],y[22]);
and and1879(ip_29_23,x[29],y[23]);
and and1880(ip_29_24,x[29],y[24]);
and and1881(ip_29_25,x[29],y[25]);
and and1882(ip_29_26,x[29],y[26]);
and and1883(ip_29_27,x[29],y[27]);
and and1884(ip_29_28,x[29],y[28]);
and and1885(ip_29_29,x[29],y[29]);
and and1886(ip_29_30,x[29],y[30]);
and and1887(ip_29_31,x[29],y[31]);
and and1888(ip_29_32,x[29],y[32]);
and and1889(ip_29_33,x[29],y[33]);
and and1890(ip_29_34,x[29],y[34]);
and and1891(ip_29_35,x[29],y[35]);
and and1892(ip_29_36,x[29],y[36]);
and and1893(ip_29_37,x[29],y[37]);
and and1894(ip_29_38,x[29],y[38]);
and and1895(ip_29_39,x[29],y[39]);
and and1896(ip_29_40,x[29],y[40]);
and and1897(ip_29_41,x[29],y[41]);
and and1898(ip_29_42,x[29],y[42]);
and and1899(ip_29_43,x[29],y[43]);
and and1900(ip_29_44,x[29],y[44]);
and and1901(ip_29_45,x[29],y[45]);
and and1902(ip_29_46,x[29],y[46]);
and and1903(ip_29_47,x[29],y[47]);
and and1904(ip_29_48,x[29],y[48]);
and and1905(ip_29_49,x[29],y[49]);
and and1906(ip_29_50,x[29],y[50]);
and and1907(ip_29_51,x[29],y[51]);
and and1908(ip_29_52,x[29],y[52]);
and and1909(ip_29_53,x[29],y[53]);
and and1910(ip_29_54,x[29],y[54]);
and and1911(ip_29_55,x[29],y[55]);
and and1912(ip_29_56,x[29],y[56]);
and and1913(ip_29_57,x[29],y[57]);
and and1914(ip_29_58,x[29],y[58]);
and and1915(ip_29_59,x[29],y[59]);
and and1916(ip_29_60,x[29],y[60]);
and and1917(ip_29_61,x[29],y[61]);
and and1918(ip_29_62,x[29],y[62]);
and and1919(ip_29_63,x[29],y[63]);
and and1920(ip_30_0,x[30],y[0]);
and and1921(ip_30_1,x[30],y[1]);
and and1922(ip_30_2,x[30],y[2]);
and and1923(ip_30_3,x[30],y[3]);
and and1924(ip_30_4,x[30],y[4]);
and and1925(ip_30_5,x[30],y[5]);
and and1926(ip_30_6,x[30],y[6]);
and and1927(ip_30_7,x[30],y[7]);
and and1928(ip_30_8,x[30],y[8]);
and and1929(ip_30_9,x[30],y[9]);
and and1930(ip_30_10,x[30],y[10]);
and and1931(ip_30_11,x[30],y[11]);
and and1932(ip_30_12,x[30],y[12]);
and and1933(ip_30_13,x[30],y[13]);
and and1934(ip_30_14,x[30],y[14]);
and and1935(ip_30_15,x[30],y[15]);
and and1936(ip_30_16,x[30],y[16]);
and and1937(ip_30_17,x[30],y[17]);
and and1938(ip_30_18,x[30],y[18]);
and and1939(ip_30_19,x[30],y[19]);
and and1940(ip_30_20,x[30],y[20]);
and and1941(ip_30_21,x[30],y[21]);
and and1942(ip_30_22,x[30],y[22]);
and and1943(ip_30_23,x[30],y[23]);
and and1944(ip_30_24,x[30],y[24]);
and and1945(ip_30_25,x[30],y[25]);
and and1946(ip_30_26,x[30],y[26]);
and and1947(ip_30_27,x[30],y[27]);
and and1948(ip_30_28,x[30],y[28]);
and and1949(ip_30_29,x[30],y[29]);
and and1950(ip_30_30,x[30],y[30]);
and and1951(ip_30_31,x[30],y[31]);
and and1952(ip_30_32,x[30],y[32]);
and and1953(ip_30_33,x[30],y[33]);
and and1954(ip_30_34,x[30],y[34]);
and and1955(ip_30_35,x[30],y[35]);
and and1956(ip_30_36,x[30],y[36]);
and and1957(ip_30_37,x[30],y[37]);
and and1958(ip_30_38,x[30],y[38]);
and and1959(ip_30_39,x[30],y[39]);
and and1960(ip_30_40,x[30],y[40]);
and and1961(ip_30_41,x[30],y[41]);
and and1962(ip_30_42,x[30],y[42]);
and and1963(ip_30_43,x[30],y[43]);
and and1964(ip_30_44,x[30],y[44]);
and and1965(ip_30_45,x[30],y[45]);
and and1966(ip_30_46,x[30],y[46]);
and and1967(ip_30_47,x[30],y[47]);
and and1968(ip_30_48,x[30],y[48]);
and and1969(ip_30_49,x[30],y[49]);
and and1970(ip_30_50,x[30],y[50]);
and and1971(ip_30_51,x[30],y[51]);
and and1972(ip_30_52,x[30],y[52]);
and and1973(ip_30_53,x[30],y[53]);
and and1974(ip_30_54,x[30],y[54]);
and and1975(ip_30_55,x[30],y[55]);
and and1976(ip_30_56,x[30],y[56]);
and and1977(ip_30_57,x[30],y[57]);
and and1978(ip_30_58,x[30],y[58]);
and and1979(ip_30_59,x[30],y[59]);
and and1980(ip_30_60,x[30],y[60]);
and and1981(ip_30_61,x[30],y[61]);
and and1982(ip_30_62,x[30],y[62]);
and and1983(ip_30_63,x[30],y[63]);
and and1984(ip_31_0,x[31],y[0]);
and and1985(ip_31_1,x[31],y[1]);
and and1986(ip_31_2,x[31],y[2]);
and and1987(ip_31_3,x[31],y[3]);
and and1988(ip_31_4,x[31],y[4]);
and and1989(ip_31_5,x[31],y[5]);
and and1990(ip_31_6,x[31],y[6]);
and and1991(ip_31_7,x[31],y[7]);
and and1992(ip_31_8,x[31],y[8]);
and and1993(ip_31_9,x[31],y[9]);
and and1994(ip_31_10,x[31],y[10]);
and and1995(ip_31_11,x[31],y[11]);
and and1996(ip_31_12,x[31],y[12]);
and and1997(ip_31_13,x[31],y[13]);
and and1998(ip_31_14,x[31],y[14]);
and and1999(ip_31_15,x[31],y[15]);
and and2000(ip_31_16,x[31],y[16]);
and and2001(ip_31_17,x[31],y[17]);
and and2002(ip_31_18,x[31],y[18]);
and and2003(ip_31_19,x[31],y[19]);
and and2004(ip_31_20,x[31],y[20]);
and and2005(ip_31_21,x[31],y[21]);
and and2006(ip_31_22,x[31],y[22]);
and and2007(ip_31_23,x[31],y[23]);
and and2008(ip_31_24,x[31],y[24]);
and and2009(ip_31_25,x[31],y[25]);
and and2010(ip_31_26,x[31],y[26]);
and and2011(ip_31_27,x[31],y[27]);
and and2012(ip_31_28,x[31],y[28]);
and and2013(ip_31_29,x[31],y[29]);
and and2014(ip_31_30,x[31],y[30]);
and and2015(ip_31_31,x[31],y[31]);
and and2016(ip_31_32,x[31],y[32]);
and and2017(ip_31_33,x[31],y[33]);
and and2018(ip_31_34,x[31],y[34]);
and and2019(ip_31_35,x[31],y[35]);
and and2020(ip_31_36,x[31],y[36]);
and and2021(ip_31_37,x[31],y[37]);
and and2022(ip_31_38,x[31],y[38]);
and and2023(ip_31_39,x[31],y[39]);
and and2024(ip_31_40,x[31],y[40]);
and and2025(ip_31_41,x[31],y[41]);
and and2026(ip_31_42,x[31],y[42]);
and and2027(ip_31_43,x[31],y[43]);
and and2028(ip_31_44,x[31],y[44]);
and and2029(ip_31_45,x[31],y[45]);
and and2030(ip_31_46,x[31],y[46]);
and and2031(ip_31_47,x[31],y[47]);
and and2032(ip_31_48,x[31],y[48]);
and and2033(ip_31_49,x[31],y[49]);
and and2034(ip_31_50,x[31],y[50]);
and and2035(ip_31_51,x[31],y[51]);
and and2036(ip_31_52,x[31],y[52]);
and and2037(ip_31_53,x[31],y[53]);
and and2038(ip_31_54,x[31],y[54]);
and and2039(ip_31_55,x[31],y[55]);
and and2040(ip_31_56,x[31],y[56]);
and and2041(ip_31_57,x[31],y[57]);
and and2042(ip_31_58,x[31],y[58]);
and and2043(ip_31_59,x[31],y[59]);
and and2044(ip_31_60,x[31],y[60]);
and and2045(ip_31_61,x[31],y[61]);
and and2046(ip_31_62,x[31],y[62]);
and and2047(ip_31_63,x[31],y[63]);
and and2048(ip_32_0,x[32],y[0]);
and and2049(ip_32_1,x[32],y[1]);
and and2050(ip_32_2,x[32],y[2]);
and and2051(ip_32_3,x[32],y[3]);
and and2052(ip_32_4,x[32],y[4]);
and and2053(ip_32_5,x[32],y[5]);
and and2054(ip_32_6,x[32],y[6]);
and and2055(ip_32_7,x[32],y[7]);
and and2056(ip_32_8,x[32],y[8]);
and and2057(ip_32_9,x[32],y[9]);
and and2058(ip_32_10,x[32],y[10]);
and and2059(ip_32_11,x[32],y[11]);
and and2060(ip_32_12,x[32],y[12]);
and and2061(ip_32_13,x[32],y[13]);
and and2062(ip_32_14,x[32],y[14]);
and and2063(ip_32_15,x[32],y[15]);
and and2064(ip_32_16,x[32],y[16]);
and and2065(ip_32_17,x[32],y[17]);
and and2066(ip_32_18,x[32],y[18]);
and and2067(ip_32_19,x[32],y[19]);
and and2068(ip_32_20,x[32],y[20]);
and and2069(ip_32_21,x[32],y[21]);
and and2070(ip_32_22,x[32],y[22]);
and and2071(ip_32_23,x[32],y[23]);
and and2072(ip_32_24,x[32],y[24]);
and and2073(ip_32_25,x[32],y[25]);
and and2074(ip_32_26,x[32],y[26]);
and and2075(ip_32_27,x[32],y[27]);
and and2076(ip_32_28,x[32],y[28]);
and and2077(ip_32_29,x[32],y[29]);
and and2078(ip_32_30,x[32],y[30]);
and and2079(ip_32_31,x[32],y[31]);
and and2080(ip_32_32,x[32],y[32]);
and and2081(ip_32_33,x[32],y[33]);
and and2082(ip_32_34,x[32],y[34]);
and and2083(ip_32_35,x[32],y[35]);
and and2084(ip_32_36,x[32],y[36]);
and and2085(ip_32_37,x[32],y[37]);
and and2086(ip_32_38,x[32],y[38]);
and and2087(ip_32_39,x[32],y[39]);
and and2088(ip_32_40,x[32],y[40]);
and and2089(ip_32_41,x[32],y[41]);
and and2090(ip_32_42,x[32],y[42]);
and and2091(ip_32_43,x[32],y[43]);
and and2092(ip_32_44,x[32],y[44]);
and and2093(ip_32_45,x[32],y[45]);
and and2094(ip_32_46,x[32],y[46]);
and and2095(ip_32_47,x[32],y[47]);
and and2096(ip_32_48,x[32],y[48]);
and and2097(ip_32_49,x[32],y[49]);
and and2098(ip_32_50,x[32],y[50]);
and and2099(ip_32_51,x[32],y[51]);
and and2100(ip_32_52,x[32],y[52]);
and and2101(ip_32_53,x[32],y[53]);
and and2102(ip_32_54,x[32],y[54]);
and and2103(ip_32_55,x[32],y[55]);
and and2104(ip_32_56,x[32],y[56]);
and and2105(ip_32_57,x[32],y[57]);
and and2106(ip_32_58,x[32],y[58]);
and and2107(ip_32_59,x[32],y[59]);
and and2108(ip_32_60,x[32],y[60]);
and and2109(ip_32_61,x[32],y[61]);
and and2110(ip_32_62,x[32],y[62]);
and and2111(ip_32_63,x[32],y[63]);
and and2112(ip_33_0,x[33],y[0]);
and and2113(ip_33_1,x[33],y[1]);
and and2114(ip_33_2,x[33],y[2]);
and and2115(ip_33_3,x[33],y[3]);
and and2116(ip_33_4,x[33],y[4]);
and and2117(ip_33_5,x[33],y[5]);
and and2118(ip_33_6,x[33],y[6]);
and and2119(ip_33_7,x[33],y[7]);
and and2120(ip_33_8,x[33],y[8]);
and and2121(ip_33_9,x[33],y[9]);
and and2122(ip_33_10,x[33],y[10]);
and and2123(ip_33_11,x[33],y[11]);
and and2124(ip_33_12,x[33],y[12]);
and and2125(ip_33_13,x[33],y[13]);
and and2126(ip_33_14,x[33],y[14]);
and and2127(ip_33_15,x[33],y[15]);
and and2128(ip_33_16,x[33],y[16]);
and and2129(ip_33_17,x[33],y[17]);
and and2130(ip_33_18,x[33],y[18]);
and and2131(ip_33_19,x[33],y[19]);
and and2132(ip_33_20,x[33],y[20]);
and and2133(ip_33_21,x[33],y[21]);
and and2134(ip_33_22,x[33],y[22]);
and and2135(ip_33_23,x[33],y[23]);
and and2136(ip_33_24,x[33],y[24]);
and and2137(ip_33_25,x[33],y[25]);
and and2138(ip_33_26,x[33],y[26]);
and and2139(ip_33_27,x[33],y[27]);
and and2140(ip_33_28,x[33],y[28]);
and and2141(ip_33_29,x[33],y[29]);
and and2142(ip_33_30,x[33],y[30]);
and and2143(ip_33_31,x[33],y[31]);
and and2144(ip_33_32,x[33],y[32]);
and and2145(ip_33_33,x[33],y[33]);
and and2146(ip_33_34,x[33],y[34]);
and and2147(ip_33_35,x[33],y[35]);
and and2148(ip_33_36,x[33],y[36]);
and and2149(ip_33_37,x[33],y[37]);
and and2150(ip_33_38,x[33],y[38]);
and and2151(ip_33_39,x[33],y[39]);
and and2152(ip_33_40,x[33],y[40]);
and and2153(ip_33_41,x[33],y[41]);
and and2154(ip_33_42,x[33],y[42]);
and and2155(ip_33_43,x[33],y[43]);
and and2156(ip_33_44,x[33],y[44]);
and and2157(ip_33_45,x[33],y[45]);
and and2158(ip_33_46,x[33],y[46]);
and and2159(ip_33_47,x[33],y[47]);
and and2160(ip_33_48,x[33],y[48]);
and and2161(ip_33_49,x[33],y[49]);
and and2162(ip_33_50,x[33],y[50]);
and and2163(ip_33_51,x[33],y[51]);
and and2164(ip_33_52,x[33],y[52]);
and and2165(ip_33_53,x[33],y[53]);
and and2166(ip_33_54,x[33],y[54]);
and and2167(ip_33_55,x[33],y[55]);
and and2168(ip_33_56,x[33],y[56]);
and and2169(ip_33_57,x[33],y[57]);
and and2170(ip_33_58,x[33],y[58]);
and and2171(ip_33_59,x[33],y[59]);
and and2172(ip_33_60,x[33],y[60]);
and and2173(ip_33_61,x[33],y[61]);
and and2174(ip_33_62,x[33],y[62]);
and and2175(ip_33_63,x[33],y[63]);
and and2176(ip_34_0,x[34],y[0]);
and and2177(ip_34_1,x[34],y[1]);
and and2178(ip_34_2,x[34],y[2]);
and and2179(ip_34_3,x[34],y[3]);
and and2180(ip_34_4,x[34],y[4]);
and and2181(ip_34_5,x[34],y[5]);
and and2182(ip_34_6,x[34],y[6]);
and and2183(ip_34_7,x[34],y[7]);
and and2184(ip_34_8,x[34],y[8]);
and and2185(ip_34_9,x[34],y[9]);
and and2186(ip_34_10,x[34],y[10]);
and and2187(ip_34_11,x[34],y[11]);
and and2188(ip_34_12,x[34],y[12]);
and and2189(ip_34_13,x[34],y[13]);
and and2190(ip_34_14,x[34],y[14]);
and and2191(ip_34_15,x[34],y[15]);
and and2192(ip_34_16,x[34],y[16]);
and and2193(ip_34_17,x[34],y[17]);
and and2194(ip_34_18,x[34],y[18]);
and and2195(ip_34_19,x[34],y[19]);
and and2196(ip_34_20,x[34],y[20]);
and and2197(ip_34_21,x[34],y[21]);
and and2198(ip_34_22,x[34],y[22]);
and and2199(ip_34_23,x[34],y[23]);
and and2200(ip_34_24,x[34],y[24]);
and and2201(ip_34_25,x[34],y[25]);
and and2202(ip_34_26,x[34],y[26]);
and and2203(ip_34_27,x[34],y[27]);
and and2204(ip_34_28,x[34],y[28]);
and and2205(ip_34_29,x[34],y[29]);
and and2206(ip_34_30,x[34],y[30]);
and and2207(ip_34_31,x[34],y[31]);
and and2208(ip_34_32,x[34],y[32]);
and and2209(ip_34_33,x[34],y[33]);
and and2210(ip_34_34,x[34],y[34]);
and and2211(ip_34_35,x[34],y[35]);
and and2212(ip_34_36,x[34],y[36]);
and and2213(ip_34_37,x[34],y[37]);
and and2214(ip_34_38,x[34],y[38]);
and and2215(ip_34_39,x[34],y[39]);
and and2216(ip_34_40,x[34],y[40]);
and and2217(ip_34_41,x[34],y[41]);
and and2218(ip_34_42,x[34],y[42]);
and and2219(ip_34_43,x[34],y[43]);
and and2220(ip_34_44,x[34],y[44]);
and and2221(ip_34_45,x[34],y[45]);
and and2222(ip_34_46,x[34],y[46]);
and and2223(ip_34_47,x[34],y[47]);
and and2224(ip_34_48,x[34],y[48]);
and and2225(ip_34_49,x[34],y[49]);
and and2226(ip_34_50,x[34],y[50]);
and and2227(ip_34_51,x[34],y[51]);
and and2228(ip_34_52,x[34],y[52]);
and and2229(ip_34_53,x[34],y[53]);
and and2230(ip_34_54,x[34],y[54]);
and and2231(ip_34_55,x[34],y[55]);
and and2232(ip_34_56,x[34],y[56]);
and and2233(ip_34_57,x[34],y[57]);
and and2234(ip_34_58,x[34],y[58]);
and and2235(ip_34_59,x[34],y[59]);
and and2236(ip_34_60,x[34],y[60]);
and and2237(ip_34_61,x[34],y[61]);
and and2238(ip_34_62,x[34],y[62]);
and and2239(ip_34_63,x[34],y[63]);
and and2240(ip_35_0,x[35],y[0]);
and and2241(ip_35_1,x[35],y[1]);
and and2242(ip_35_2,x[35],y[2]);
and and2243(ip_35_3,x[35],y[3]);
and and2244(ip_35_4,x[35],y[4]);
and and2245(ip_35_5,x[35],y[5]);
and and2246(ip_35_6,x[35],y[6]);
and and2247(ip_35_7,x[35],y[7]);
and and2248(ip_35_8,x[35],y[8]);
and and2249(ip_35_9,x[35],y[9]);
and and2250(ip_35_10,x[35],y[10]);
and and2251(ip_35_11,x[35],y[11]);
and and2252(ip_35_12,x[35],y[12]);
and and2253(ip_35_13,x[35],y[13]);
and and2254(ip_35_14,x[35],y[14]);
and and2255(ip_35_15,x[35],y[15]);
and and2256(ip_35_16,x[35],y[16]);
and and2257(ip_35_17,x[35],y[17]);
and and2258(ip_35_18,x[35],y[18]);
and and2259(ip_35_19,x[35],y[19]);
and and2260(ip_35_20,x[35],y[20]);
and and2261(ip_35_21,x[35],y[21]);
and and2262(ip_35_22,x[35],y[22]);
and and2263(ip_35_23,x[35],y[23]);
and and2264(ip_35_24,x[35],y[24]);
and and2265(ip_35_25,x[35],y[25]);
and and2266(ip_35_26,x[35],y[26]);
and and2267(ip_35_27,x[35],y[27]);
and and2268(ip_35_28,x[35],y[28]);
and and2269(ip_35_29,x[35],y[29]);
and and2270(ip_35_30,x[35],y[30]);
and and2271(ip_35_31,x[35],y[31]);
and and2272(ip_35_32,x[35],y[32]);
and and2273(ip_35_33,x[35],y[33]);
and and2274(ip_35_34,x[35],y[34]);
and and2275(ip_35_35,x[35],y[35]);
and and2276(ip_35_36,x[35],y[36]);
and and2277(ip_35_37,x[35],y[37]);
and and2278(ip_35_38,x[35],y[38]);
and and2279(ip_35_39,x[35],y[39]);
and and2280(ip_35_40,x[35],y[40]);
and and2281(ip_35_41,x[35],y[41]);
and and2282(ip_35_42,x[35],y[42]);
and and2283(ip_35_43,x[35],y[43]);
and and2284(ip_35_44,x[35],y[44]);
and and2285(ip_35_45,x[35],y[45]);
and and2286(ip_35_46,x[35],y[46]);
and and2287(ip_35_47,x[35],y[47]);
and and2288(ip_35_48,x[35],y[48]);
and and2289(ip_35_49,x[35],y[49]);
and and2290(ip_35_50,x[35],y[50]);
and and2291(ip_35_51,x[35],y[51]);
and and2292(ip_35_52,x[35],y[52]);
and and2293(ip_35_53,x[35],y[53]);
and and2294(ip_35_54,x[35],y[54]);
and and2295(ip_35_55,x[35],y[55]);
and and2296(ip_35_56,x[35],y[56]);
and and2297(ip_35_57,x[35],y[57]);
and and2298(ip_35_58,x[35],y[58]);
and and2299(ip_35_59,x[35],y[59]);
and and2300(ip_35_60,x[35],y[60]);
and and2301(ip_35_61,x[35],y[61]);
and and2302(ip_35_62,x[35],y[62]);
and and2303(ip_35_63,x[35],y[63]);
and and2304(ip_36_0,x[36],y[0]);
and and2305(ip_36_1,x[36],y[1]);
and and2306(ip_36_2,x[36],y[2]);
and and2307(ip_36_3,x[36],y[3]);
and and2308(ip_36_4,x[36],y[4]);
and and2309(ip_36_5,x[36],y[5]);
and and2310(ip_36_6,x[36],y[6]);
and and2311(ip_36_7,x[36],y[7]);
and and2312(ip_36_8,x[36],y[8]);
and and2313(ip_36_9,x[36],y[9]);
and and2314(ip_36_10,x[36],y[10]);
and and2315(ip_36_11,x[36],y[11]);
and and2316(ip_36_12,x[36],y[12]);
and and2317(ip_36_13,x[36],y[13]);
and and2318(ip_36_14,x[36],y[14]);
and and2319(ip_36_15,x[36],y[15]);
and and2320(ip_36_16,x[36],y[16]);
and and2321(ip_36_17,x[36],y[17]);
and and2322(ip_36_18,x[36],y[18]);
and and2323(ip_36_19,x[36],y[19]);
and and2324(ip_36_20,x[36],y[20]);
and and2325(ip_36_21,x[36],y[21]);
and and2326(ip_36_22,x[36],y[22]);
and and2327(ip_36_23,x[36],y[23]);
and and2328(ip_36_24,x[36],y[24]);
and and2329(ip_36_25,x[36],y[25]);
and and2330(ip_36_26,x[36],y[26]);
and and2331(ip_36_27,x[36],y[27]);
and and2332(ip_36_28,x[36],y[28]);
and and2333(ip_36_29,x[36],y[29]);
and and2334(ip_36_30,x[36],y[30]);
and and2335(ip_36_31,x[36],y[31]);
and and2336(ip_36_32,x[36],y[32]);
and and2337(ip_36_33,x[36],y[33]);
and and2338(ip_36_34,x[36],y[34]);
and and2339(ip_36_35,x[36],y[35]);
and and2340(ip_36_36,x[36],y[36]);
and and2341(ip_36_37,x[36],y[37]);
and and2342(ip_36_38,x[36],y[38]);
and and2343(ip_36_39,x[36],y[39]);
and and2344(ip_36_40,x[36],y[40]);
and and2345(ip_36_41,x[36],y[41]);
and and2346(ip_36_42,x[36],y[42]);
and and2347(ip_36_43,x[36],y[43]);
and and2348(ip_36_44,x[36],y[44]);
and and2349(ip_36_45,x[36],y[45]);
and and2350(ip_36_46,x[36],y[46]);
and and2351(ip_36_47,x[36],y[47]);
and and2352(ip_36_48,x[36],y[48]);
and and2353(ip_36_49,x[36],y[49]);
and and2354(ip_36_50,x[36],y[50]);
and and2355(ip_36_51,x[36],y[51]);
and and2356(ip_36_52,x[36],y[52]);
and and2357(ip_36_53,x[36],y[53]);
and and2358(ip_36_54,x[36],y[54]);
and and2359(ip_36_55,x[36],y[55]);
and and2360(ip_36_56,x[36],y[56]);
and and2361(ip_36_57,x[36],y[57]);
and and2362(ip_36_58,x[36],y[58]);
and and2363(ip_36_59,x[36],y[59]);
and and2364(ip_36_60,x[36],y[60]);
and and2365(ip_36_61,x[36],y[61]);
and and2366(ip_36_62,x[36],y[62]);
and and2367(ip_36_63,x[36],y[63]);
and and2368(ip_37_0,x[37],y[0]);
and and2369(ip_37_1,x[37],y[1]);
and and2370(ip_37_2,x[37],y[2]);
and and2371(ip_37_3,x[37],y[3]);
and and2372(ip_37_4,x[37],y[4]);
and and2373(ip_37_5,x[37],y[5]);
and and2374(ip_37_6,x[37],y[6]);
and and2375(ip_37_7,x[37],y[7]);
and and2376(ip_37_8,x[37],y[8]);
and and2377(ip_37_9,x[37],y[9]);
and and2378(ip_37_10,x[37],y[10]);
and and2379(ip_37_11,x[37],y[11]);
and and2380(ip_37_12,x[37],y[12]);
and and2381(ip_37_13,x[37],y[13]);
and and2382(ip_37_14,x[37],y[14]);
and and2383(ip_37_15,x[37],y[15]);
and and2384(ip_37_16,x[37],y[16]);
and and2385(ip_37_17,x[37],y[17]);
and and2386(ip_37_18,x[37],y[18]);
and and2387(ip_37_19,x[37],y[19]);
and and2388(ip_37_20,x[37],y[20]);
and and2389(ip_37_21,x[37],y[21]);
and and2390(ip_37_22,x[37],y[22]);
and and2391(ip_37_23,x[37],y[23]);
and and2392(ip_37_24,x[37],y[24]);
and and2393(ip_37_25,x[37],y[25]);
and and2394(ip_37_26,x[37],y[26]);
and and2395(ip_37_27,x[37],y[27]);
and and2396(ip_37_28,x[37],y[28]);
and and2397(ip_37_29,x[37],y[29]);
and and2398(ip_37_30,x[37],y[30]);
and and2399(ip_37_31,x[37],y[31]);
and and2400(ip_37_32,x[37],y[32]);
and and2401(ip_37_33,x[37],y[33]);
and and2402(ip_37_34,x[37],y[34]);
and and2403(ip_37_35,x[37],y[35]);
and and2404(ip_37_36,x[37],y[36]);
and and2405(ip_37_37,x[37],y[37]);
and and2406(ip_37_38,x[37],y[38]);
and and2407(ip_37_39,x[37],y[39]);
and and2408(ip_37_40,x[37],y[40]);
and and2409(ip_37_41,x[37],y[41]);
and and2410(ip_37_42,x[37],y[42]);
and and2411(ip_37_43,x[37],y[43]);
and and2412(ip_37_44,x[37],y[44]);
and and2413(ip_37_45,x[37],y[45]);
and and2414(ip_37_46,x[37],y[46]);
and and2415(ip_37_47,x[37],y[47]);
and and2416(ip_37_48,x[37],y[48]);
and and2417(ip_37_49,x[37],y[49]);
and and2418(ip_37_50,x[37],y[50]);
and and2419(ip_37_51,x[37],y[51]);
and and2420(ip_37_52,x[37],y[52]);
and and2421(ip_37_53,x[37],y[53]);
and and2422(ip_37_54,x[37],y[54]);
and and2423(ip_37_55,x[37],y[55]);
and and2424(ip_37_56,x[37],y[56]);
and and2425(ip_37_57,x[37],y[57]);
and and2426(ip_37_58,x[37],y[58]);
and and2427(ip_37_59,x[37],y[59]);
and and2428(ip_37_60,x[37],y[60]);
and and2429(ip_37_61,x[37],y[61]);
and and2430(ip_37_62,x[37],y[62]);
and and2431(ip_37_63,x[37],y[63]);
and and2432(ip_38_0,x[38],y[0]);
and and2433(ip_38_1,x[38],y[1]);
and and2434(ip_38_2,x[38],y[2]);
and and2435(ip_38_3,x[38],y[3]);
and and2436(ip_38_4,x[38],y[4]);
and and2437(ip_38_5,x[38],y[5]);
and and2438(ip_38_6,x[38],y[6]);
and and2439(ip_38_7,x[38],y[7]);
and and2440(ip_38_8,x[38],y[8]);
and and2441(ip_38_9,x[38],y[9]);
and and2442(ip_38_10,x[38],y[10]);
and and2443(ip_38_11,x[38],y[11]);
and and2444(ip_38_12,x[38],y[12]);
and and2445(ip_38_13,x[38],y[13]);
and and2446(ip_38_14,x[38],y[14]);
and and2447(ip_38_15,x[38],y[15]);
and and2448(ip_38_16,x[38],y[16]);
and and2449(ip_38_17,x[38],y[17]);
and and2450(ip_38_18,x[38],y[18]);
and and2451(ip_38_19,x[38],y[19]);
and and2452(ip_38_20,x[38],y[20]);
and and2453(ip_38_21,x[38],y[21]);
and and2454(ip_38_22,x[38],y[22]);
and and2455(ip_38_23,x[38],y[23]);
and and2456(ip_38_24,x[38],y[24]);
and and2457(ip_38_25,x[38],y[25]);
and and2458(ip_38_26,x[38],y[26]);
and and2459(ip_38_27,x[38],y[27]);
and and2460(ip_38_28,x[38],y[28]);
and and2461(ip_38_29,x[38],y[29]);
and and2462(ip_38_30,x[38],y[30]);
and and2463(ip_38_31,x[38],y[31]);
and and2464(ip_38_32,x[38],y[32]);
and and2465(ip_38_33,x[38],y[33]);
and and2466(ip_38_34,x[38],y[34]);
and and2467(ip_38_35,x[38],y[35]);
and and2468(ip_38_36,x[38],y[36]);
and and2469(ip_38_37,x[38],y[37]);
and and2470(ip_38_38,x[38],y[38]);
and and2471(ip_38_39,x[38],y[39]);
and and2472(ip_38_40,x[38],y[40]);
and and2473(ip_38_41,x[38],y[41]);
and and2474(ip_38_42,x[38],y[42]);
and and2475(ip_38_43,x[38],y[43]);
and and2476(ip_38_44,x[38],y[44]);
and and2477(ip_38_45,x[38],y[45]);
and and2478(ip_38_46,x[38],y[46]);
and and2479(ip_38_47,x[38],y[47]);
and and2480(ip_38_48,x[38],y[48]);
and and2481(ip_38_49,x[38],y[49]);
and and2482(ip_38_50,x[38],y[50]);
and and2483(ip_38_51,x[38],y[51]);
and and2484(ip_38_52,x[38],y[52]);
and and2485(ip_38_53,x[38],y[53]);
and and2486(ip_38_54,x[38],y[54]);
and and2487(ip_38_55,x[38],y[55]);
and and2488(ip_38_56,x[38],y[56]);
and and2489(ip_38_57,x[38],y[57]);
and and2490(ip_38_58,x[38],y[58]);
and and2491(ip_38_59,x[38],y[59]);
and and2492(ip_38_60,x[38],y[60]);
and and2493(ip_38_61,x[38],y[61]);
and and2494(ip_38_62,x[38],y[62]);
and and2495(ip_38_63,x[38],y[63]);
and and2496(ip_39_0,x[39],y[0]);
and and2497(ip_39_1,x[39],y[1]);
and and2498(ip_39_2,x[39],y[2]);
and and2499(ip_39_3,x[39],y[3]);
and and2500(ip_39_4,x[39],y[4]);
and and2501(ip_39_5,x[39],y[5]);
and and2502(ip_39_6,x[39],y[6]);
and and2503(ip_39_7,x[39],y[7]);
and and2504(ip_39_8,x[39],y[8]);
and and2505(ip_39_9,x[39],y[9]);
and and2506(ip_39_10,x[39],y[10]);
and and2507(ip_39_11,x[39],y[11]);
and and2508(ip_39_12,x[39],y[12]);
and and2509(ip_39_13,x[39],y[13]);
and and2510(ip_39_14,x[39],y[14]);
and and2511(ip_39_15,x[39],y[15]);
and and2512(ip_39_16,x[39],y[16]);
and and2513(ip_39_17,x[39],y[17]);
and and2514(ip_39_18,x[39],y[18]);
and and2515(ip_39_19,x[39],y[19]);
and and2516(ip_39_20,x[39],y[20]);
and and2517(ip_39_21,x[39],y[21]);
and and2518(ip_39_22,x[39],y[22]);
and and2519(ip_39_23,x[39],y[23]);
and and2520(ip_39_24,x[39],y[24]);
and and2521(ip_39_25,x[39],y[25]);
and and2522(ip_39_26,x[39],y[26]);
and and2523(ip_39_27,x[39],y[27]);
and and2524(ip_39_28,x[39],y[28]);
and and2525(ip_39_29,x[39],y[29]);
and and2526(ip_39_30,x[39],y[30]);
and and2527(ip_39_31,x[39],y[31]);
and and2528(ip_39_32,x[39],y[32]);
and and2529(ip_39_33,x[39],y[33]);
and and2530(ip_39_34,x[39],y[34]);
and and2531(ip_39_35,x[39],y[35]);
and and2532(ip_39_36,x[39],y[36]);
and and2533(ip_39_37,x[39],y[37]);
and and2534(ip_39_38,x[39],y[38]);
and and2535(ip_39_39,x[39],y[39]);
and and2536(ip_39_40,x[39],y[40]);
and and2537(ip_39_41,x[39],y[41]);
and and2538(ip_39_42,x[39],y[42]);
and and2539(ip_39_43,x[39],y[43]);
and and2540(ip_39_44,x[39],y[44]);
and and2541(ip_39_45,x[39],y[45]);
and and2542(ip_39_46,x[39],y[46]);
and and2543(ip_39_47,x[39],y[47]);
and and2544(ip_39_48,x[39],y[48]);
and and2545(ip_39_49,x[39],y[49]);
and and2546(ip_39_50,x[39],y[50]);
and and2547(ip_39_51,x[39],y[51]);
and and2548(ip_39_52,x[39],y[52]);
and and2549(ip_39_53,x[39],y[53]);
and and2550(ip_39_54,x[39],y[54]);
and and2551(ip_39_55,x[39],y[55]);
and and2552(ip_39_56,x[39],y[56]);
and and2553(ip_39_57,x[39],y[57]);
and and2554(ip_39_58,x[39],y[58]);
and and2555(ip_39_59,x[39],y[59]);
and and2556(ip_39_60,x[39],y[60]);
and and2557(ip_39_61,x[39],y[61]);
and and2558(ip_39_62,x[39],y[62]);
and and2559(ip_39_63,x[39],y[63]);
and and2560(ip_40_0,x[40],y[0]);
and and2561(ip_40_1,x[40],y[1]);
and and2562(ip_40_2,x[40],y[2]);
and and2563(ip_40_3,x[40],y[3]);
and and2564(ip_40_4,x[40],y[4]);
and and2565(ip_40_5,x[40],y[5]);
and and2566(ip_40_6,x[40],y[6]);
and and2567(ip_40_7,x[40],y[7]);
and and2568(ip_40_8,x[40],y[8]);
and and2569(ip_40_9,x[40],y[9]);
and and2570(ip_40_10,x[40],y[10]);
and and2571(ip_40_11,x[40],y[11]);
and and2572(ip_40_12,x[40],y[12]);
and and2573(ip_40_13,x[40],y[13]);
and and2574(ip_40_14,x[40],y[14]);
and and2575(ip_40_15,x[40],y[15]);
and and2576(ip_40_16,x[40],y[16]);
and and2577(ip_40_17,x[40],y[17]);
and and2578(ip_40_18,x[40],y[18]);
and and2579(ip_40_19,x[40],y[19]);
and and2580(ip_40_20,x[40],y[20]);
and and2581(ip_40_21,x[40],y[21]);
and and2582(ip_40_22,x[40],y[22]);
and and2583(ip_40_23,x[40],y[23]);
and and2584(ip_40_24,x[40],y[24]);
and and2585(ip_40_25,x[40],y[25]);
and and2586(ip_40_26,x[40],y[26]);
and and2587(ip_40_27,x[40],y[27]);
and and2588(ip_40_28,x[40],y[28]);
and and2589(ip_40_29,x[40],y[29]);
and and2590(ip_40_30,x[40],y[30]);
and and2591(ip_40_31,x[40],y[31]);
and and2592(ip_40_32,x[40],y[32]);
and and2593(ip_40_33,x[40],y[33]);
and and2594(ip_40_34,x[40],y[34]);
and and2595(ip_40_35,x[40],y[35]);
and and2596(ip_40_36,x[40],y[36]);
and and2597(ip_40_37,x[40],y[37]);
and and2598(ip_40_38,x[40],y[38]);
and and2599(ip_40_39,x[40],y[39]);
and and2600(ip_40_40,x[40],y[40]);
and and2601(ip_40_41,x[40],y[41]);
and and2602(ip_40_42,x[40],y[42]);
and and2603(ip_40_43,x[40],y[43]);
and and2604(ip_40_44,x[40],y[44]);
and and2605(ip_40_45,x[40],y[45]);
and and2606(ip_40_46,x[40],y[46]);
and and2607(ip_40_47,x[40],y[47]);
and and2608(ip_40_48,x[40],y[48]);
and and2609(ip_40_49,x[40],y[49]);
and and2610(ip_40_50,x[40],y[50]);
and and2611(ip_40_51,x[40],y[51]);
and and2612(ip_40_52,x[40],y[52]);
and and2613(ip_40_53,x[40],y[53]);
and and2614(ip_40_54,x[40],y[54]);
and and2615(ip_40_55,x[40],y[55]);
and and2616(ip_40_56,x[40],y[56]);
and and2617(ip_40_57,x[40],y[57]);
and and2618(ip_40_58,x[40],y[58]);
and and2619(ip_40_59,x[40],y[59]);
and and2620(ip_40_60,x[40],y[60]);
and and2621(ip_40_61,x[40],y[61]);
and and2622(ip_40_62,x[40],y[62]);
and and2623(ip_40_63,x[40],y[63]);
and and2624(ip_41_0,x[41],y[0]);
and and2625(ip_41_1,x[41],y[1]);
and and2626(ip_41_2,x[41],y[2]);
and and2627(ip_41_3,x[41],y[3]);
and and2628(ip_41_4,x[41],y[4]);
and and2629(ip_41_5,x[41],y[5]);
and and2630(ip_41_6,x[41],y[6]);
and and2631(ip_41_7,x[41],y[7]);
and and2632(ip_41_8,x[41],y[8]);
and and2633(ip_41_9,x[41],y[9]);
and and2634(ip_41_10,x[41],y[10]);
and and2635(ip_41_11,x[41],y[11]);
and and2636(ip_41_12,x[41],y[12]);
and and2637(ip_41_13,x[41],y[13]);
and and2638(ip_41_14,x[41],y[14]);
and and2639(ip_41_15,x[41],y[15]);
and and2640(ip_41_16,x[41],y[16]);
and and2641(ip_41_17,x[41],y[17]);
and and2642(ip_41_18,x[41],y[18]);
and and2643(ip_41_19,x[41],y[19]);
and and2644(ip_41_20,x[41],y[20]);
and and2645(ip_41_21,x[41],y[21]);
and and2646(ip_41_22,x[41],y[22]);
and and2647(ip_41_23,x[41],y[23]);
and and2648(ip_41_24,x[41],y[24]);
and and2649(ip_41_25,x[41],y[25]);
and and2650(ip_41_26,x[41],y[26]);
and and2651(ip_41_27,x[41],y[27]);
and and2652(ip_41_28,x[41],y[28]);
and and2653(ip_41_29,x[41],y[29]);
and and2654(ip_41_30,x[41],y[30]);
and and2655(ip_41_31,x[41],y[31]);
and and2656(ip_41_32,x[41],y[32]);
and and2657(ip_41_33,x[41],y[33]);
and and2658(ip_41_34,x[41],y[34]);
and and2659(ip_41_35,x[41],y[35]);
and and2660(ip_41_36,x[41],y[36]);
and and2661(ip_41_37,x[41],y[37]);
and and2662(ip_41_38,x[41],y[38]);
and and2663(ip_41_39,x[41],y[39]);
and and2664(ip_41_40,x[41],y[40]);
and and2665(ip_41_41,x[41],y[41]);
and and2666(ip_41_42,x[41],y[42]);
and and2667(ip_41_43,x[41],y[43]);
and and2668(ip_41_44,x[41],y[44]);
and and2669(ip_41_45,x[41],y[45]);
and and2670(ip_41_46,x[41],y[46]);
and and2671(ip_41_47,x[41],y[47]);
and and2672(ip_41_48,x[41],y[48]);
and and2673(ip_41_49,x[41],y[49]);
and and2674(ip_41_50,x[41],y[50]);
and and2675(ip_41_51,x[41],y[51]);
and and2676(ip_41_52,x[41],y[52]);
and and2677(ip_41_53,x[41],y[53]);
and and2678(ip_41_54,x[41],y[54]);
and and2679(ip_41_55,x[41],y[55]);
and and2680(ip_41_56,x[41],y[56]);
and and2681(ip_41_57,x[41],y[57]);
and and2682(ip_41_58,x[41],y[58]);
and and2683(ip_41_59,x[41],y[59]);
and and2684(ip_41_60,x[41],y[60]);
and and2685(ip_41_61,x[41],y[61]);
and and2686(ip_41_62,x[41],y[62]);
and and2687(ip_41_63,x[41],y[63]);
and and2688(ip_42_0,x[42],y[0]);
and and2689(ip_42_1,x[42],y[1]);
and and2690(ip_42_2,x[42],y[2]);
and and2691(ip_42_3,x[42],y[3]);
and and2692(ip_42_4,x[42],y[4]);
and and2693(ip_42_5,x[42],y[5]);
and and2694(ip_42_6,x[42],y[6]);
and and2695(ip_42_7,x[42],y[7]);
and and2696(ip_42_8,x[42],y[8]);
and and2697(ip_42_9,x[42],y[9]);
and and2698(ip_42_10,x[42],y[10]);
and and2699(ip_42_11,x[42],y[11]);
and and2700(ip_42_12,x[42],y[12]);
and and2701(ip_42_13,x[42],y[13]);
and and2702(ip_42_14,x[42],y[14]);
and and2703(ip_42_15,x[42],y[15]);
and and2704(ip_42_16,x[42],y[16]);
and and2705(ip_42_17,x[42],y[17]);
and and2706(ip_42_18,x[42],y[18]);
and and2707(ip_42_19,x[42],y[19]);
and and2708(ip_42_20,x[42],y[20]);
and and2709(ip_42_21,x[42],y[21]);
and and2710(ip_42_22,x[42],y[22]);
and and2711(ip_42_23,x[42],y[23]);
and and2712(ip_42_24,x[42],y[24]);
and and2713(ip_42_25,x[42],y[25]);
and and2714(ip_42_26,x[42],y[26]);
and and2715(ip_42_27,x[42],y[27]);
and and2716(ip_42_28,x[42],y[28]);
and and2717(ip_42_29,x[42],y[29]);
and and2718(ip_42_30,x[42],y[30]);
and and2719(ip_42_31,x[42],y[31]);
and and2720(ip_42_32,x[42],y[32]);
and and2721(ip_42_33,x[42],y[33]);
and and2722(ip_42_34,x[42],y[34]);
and and2723(ip_42_35,x[42],y[35]);
and and2724(ip_42_36,x[42],y[36]);
and and2725(ip_42_37,x[42],y[37]);
and and2726(ip_42_38,x[42],y[38]);
and and2727(ip_42_39,x[42],y[39]);
and and2728(ip_42_40,x[42],y[40]);
and and2729(ip_42_41,x[42],y[41]);
and and2730(ip_42_42,x[42],y[42]);
and and2731(ip_42_43,x[42],y[43]);
and and2732(ip_42_44,x[42],y[44]);
and and2733(ip_42_45,x[42],y[45]);
and and2734(ip_42_46,x[42],y[46]);
and and2735(ip_42_47,x[42],y[47]);
and and2736(ip_42_48,x[42],y[48]);
and and2737(ip_42_49,x[42],y[49]);
and and2738(ip_42_50,x[42],y[50]);
and and2739(ip_42_51,x[42],y[51]);
and and2740(ip_42_52,x[42],y[52]);
and and2741(ip_42_53,x[42],y[53]);
and and2742(ip_42_54,x[42],y[54]);
and and2743(ip_42_55,x[42],y[55]);
and and2744(ip_42_56,x[42],y[56]);
and and2745(ip_42_57,x[42],y[57]);
and and2746(ip_42_58,x[42],y[58]);
and and2747(ip_42_59,x[42],y[59]);
and and2748(ip_42_60,x[42],y[60]);
and and2749(ip_42_61,x[42],y[61]);
and and2750(ip_42_62,x[42],y[62]);
and and2751(ip_42_63,x[42],y[63]);
and and2752(ip_43_0,x[43],y[0]);
and and2753(ip_43_1,x[43],y[1]);
and and2754(ip_43_2,x[43],y[2]);
and and2755(ip_43_3,x[43],y[3]);
and and2756(ip_43_4,x[43],y[4]);
and and2757(ip_43_5,x[43],y[5]);
and and2758(ip_43_6,x[43],y[6]);
and and2759(ip_43_7,x[43],y[7]);
and and2760(ip_43_8,x[43],y[8]);
and and2761(ip_43_9,x[43],y[9]);
and and2762(ip_43_10,x[43],y[10]);
and and2763(ip_43_11,x[43],y[11]);
and and2764(ip_43_12,x[43],y[12]);
and and2765(ip_43_13,x[43],y[13]);
and and2766(ip_43_14,x[43],y[14]);
and and2767(ip_43_15,x[43],y[15]);
and and2768(ip_43_16,x[43],y[16]);
and and2769(ip_43_17,x[43],y[17]);
and and2770(ip_43_18,x[43],y[18]);
and and2771(ip_43_19,x[43],y[19]);
and and2772(ip_43_20,x[43],y[20]);
and and2773(ip_43_21,x[43],y[21]);
and and2774(ip_43_22,x[43],y[22]);
and and2775(ip_43_23,x[43],y[23]);
and and2776(ip_43_24,x[43],y[24]);
and and2777(ip_43_25,x[43],y[25]);
and and2778(ip_43_26,x[43],y[26]);
and and2779(ip_43_27,x[43],y[27]);
and and2780(ip_43_28,x[43],y[28]);
and and2781(ip_43_29,x[43],y[29]);
and and2782(ip_43_30,x[43],y[30]);
and and2783(ip_43_31,x[43],y[31]);
and and2784(ip_43_32,x[43],y[32]);
and and2785(ip_43_33,x[43],y[33]);
and and2786(ip_43_34,x[43],y[34]);
and and2787(ip_43_35,x[43],y[35]);
and and2788(ip_43_36,x[43],y[36]);
and and2789(ip_43_37,x[43],y[37]);
and and2790(ip_43_38,x[43],y[38]);
and and2791(ip_43_39,x[43],y[39]);
and and2792(ip_43_40,x[43],y[40]);
and and2793(ip_43_41,x[43],y[41]);
and and2794(ip_43_42,x[43],y[42]);
and and2795(ip_43_43,x[43],y[43]);
and and2796(ip_43_44,x[43],y[44]);
and and2797(ip_43_45,x[43],y[45]);
and and2798(ip_43_46,x[43],y[46]);
and and2799(ip_43_47,x[43],y[47]);
and and2800(ip_43_48,x[43],y[48]);
and and2801(ip_43_49,x[43],y[49]);
and and2802(ip_43_50,x[43],y[50]);
and and2803(ip_43_51,x[43],y[51]);
and and2804(ip_43_52,x[43],y[52]);
and and2805(ip_43_53,x[43],y[53]);
and and2806(ip_43_54,x[43],y[54]);
and and2807(ip_43_55,x[43],y[55]);
and and2808(ip_43_56,x[43],y[56]);
and and2809(ip_43_57,x[43],y[57]);
and and2810(ip_43_58,x[43],y[58]);
and and2811(ip_43_59,x[43],y[59]);
and and2812(ip_43_60,x[43],y[60]);
and and2813(ip_43_61,x[43],y[61]);
and and2814(ip_43_62,x[43],y[62]);
and and2815(ip_43_63,x[43],y[63]);
and and2816(ip_44_0,x[44],y[0]);
and and2817(ip_44_1,x[44],y[1]);
and and2818(ip_44_2,x[44],y[2]);
and and2819(ip_44_3,x[44],y[3]);
and and2820(ip_44_4,x[44],y[4]);
and and2821(ip_44_5,x[44],y[5]);
and and2822(ip_44_6,x[44],y[6]);
and and2823(ip_44_7,x[44],y[7]);
and and2824(ip_44_8,x[44],y[8]);
and and2825(ip_44_9,x[44],y[9]);
and and2826(ip_44_10,x[44],y[10]);
and and2827(ip_44_11,x[44],y[11]);
and and2828(ip_44_12,x[44],y[12]);
and and2829(ip_44_13,x[44],y[13]);
and and2830(ip_44_14,x[44],y[14]);
and and2831(ip_44_15,x[44],y[15]);
and and2832(ip_44_16,x[44],y[16]);
and and2833(ip_44_17,x[44],y[17]);
and and2834(ip_44_18,x[44],y[18]);
and and2835(ip_44_19,x[44],y[19]);
and and2836(ip_44_20,x[44],y[20]);
and and2837(ip_44_21,x[44],y[21]);
and and2838(ip_44_22,x[44],y[22]);
and and2839(ip_44_23,x[44],y[23]);
and and2840(ip_44_24,x[44],y[24]);
and and2841(ip_44_25,x[44],y[25]);
and and2842(ip_44_26,x[44],y[26]);
and and2843(ip_44_27,x[44],y[27]);
and and2844(ip_44_28,x[44],y[28]);
and and2845(ip_44_29,x[44],y[29]);
and and2846(ip_44_30,x[44],y[30]);
and and2847(ip_44_31,x[44],y[31]);
and and2848(ip_44_32,x[44],y[32]);
and and2849(ip_44_33,x[44],y[33]);
and and2850(ip_44_34,x[44],y[34]);
and and2851(ip_44_35,x[44],y[35]);
and and2852(ip_44_36,x[44],y[36]);
and and2853(ip_44_37,x[44],y[37]);
and and2854(ip_44_38,x[44],y[38]);
and and2855(ip_44_39,x[44],y[39]);
and and2856(ip_44_40,x[44],y[40]);
and and2857(ip_44_41,x[44],y[41]);
and and2858(ip_44_42,x[44],y[42]);
and and2859(ip_44_43,x[44],y[43]);
and and2860(ip_44_44,x[44],y[44]);
and and2861(ip_44_45,x[44],y[45]);
and and2862(ip_44_46,x[44],y[46]);
and and2863(ip_44_47,x[44],y[47]);
and and2864(ip_44_48,x[44],y[48]);
and and2865(ip_44_49,x[44],y[49]);
and and2866(ip_44_50,x[44],y[50]);
and and2867(ip_44_51,x[44],y[51]);
and and2868(ip_44_52,x[44],y[52]);
and and2869(ip_44_53,x[44],y[53]);
and and2870(ip_44_54,x[44],y[54]);
and and2871(ip_44_55,x[44],y[55]);
and and2872(ip_44_56,x[44],y[56]);
and and2873(ip_44_57,x[44],y[57]);
and and2874(ip_44_58,x[44],y[58]);
and and2875(ip_44_59,x[44],y[59]);
and and2876(ip_44_60,x[44],y[60]);
and and2877(ip_44_61,x[44],y[61]);
and and2878(ip_44_62,x[44],y[62]);
and and2879(ip_44_63,x[44],y[63]);
and and2880(ip_45_0,x[45],y[0]);
and and2881(ip_45_1,x[45],y[1]);
and and2882(ip_45_2,x[45],y[2]);
and and2883(ip_45_3,x[45],y[3]);
and and2884(ip_45_4,x[45],y[4]);
and and2885(ip_45_5,x[45],y[5]);
and and2886(ip_45_6,x[45],y[6]);
and and2887(ip_45_7,x[45],y[7]);
and and2888(ip_45_8,x[45],y[8]);
and and2889(ip_45_9,x[45],y[9]);
and and2890(ip_45_10,x[45],y[10]);
and and2891(ip_45_11,x[45],y[11]);
and and2892(ip_45_12,x[45],y[12]);
and and2893(ip_45_13,x[45],y[13]);
and and2894(ip_45_14,x[45],y[14]);
and and2895(ip_45_15,x[45],y[15]);
and and2896(ip_45_16,x[45],y[16]);
and and2897(ip_45_17,x[45],y[17]);
and and2898(ip_45_18,x[45],y[18]);
and and2899(ip_45_19,x[45],y[19]);
and and2900(ip_45_20,x[45],y[20]);
and and2901(ip_45_21,x[45],y[21]);
and and2902(ip_45_22,x[45],y[22]);
and and2903(ip_45_23,x[45],y[23]);
and and2904(ip_45_24,x[45],y[24]);
and and2905(ip_45_25,x[45],y[25]);
and and2906(ip_45_26,x[45],y[26]);
and and2907(ip_45_27,x[45],y[27]);
and and2908(ip_45_28,x[45],y[28]);
and and2909(ip_45_29,x[45],y[29]);
and and2910(ip_45_30,x[45],y[30]);
and and2911(ip_45_31,x[45],y[31]);
and and2912(ip_45_32,x[45],y[32]);
and and2913(ip_45_33,x[45],y[33]);
and and2914(ip_45_34,x[45],y[34]);
and and2915(ip_45_35,x[45],y[35]);
and and2916(ip_45_36,x[45],y[36]);
and and2917(ip_45_37,x[45],y[37]);
and and2918(ip_45_38,x[45],y[38]);
and and2919(ip_45_39,x[45],y[39]);
and and2920(ip_45_40,x[45],y[40]);
and and2921(ip_45_41,x[45],y[41]);
and and2922(ip_45_42,x[45],y[42]);
and and2923(ip_45_43,x[45],y[43]);
and and2924(ip_45_44,x[45],y[44]);
and and2925(ip_45_45,x[45],y[45]);
and and2926(ip_45_46,x[45],y[46]);
and and2927(ip_45_47,x[45],y[47]);
and and2928(ip_45_48,x[45],y[48]);
and and2929(ip_45_49,x[45],y[49]);
and and2930(ip_45_50,x[45],y[50]);
and and2931(ip_45_51,x[45],y[51]);
and and2932(ip_45_52,x[45],y[52]);
and and2933(ip_45_53,x[45],y[53]);
and and2934(ip_45_54,x[45],y[54]);
and and2935(ip_45_55,x[45],y[55]);
and and2936(ip_45_56,x[45],y[56]);
and and2937(ip_45_57,x[45],y[57]);
and and2938(ip_45_58,x[45],y[58]);
and and2939(ip_45_59,x[45],y[59]);
and and2940(ip_45_60,x[45],y[60]);
and and2941(ip_45_61,x[45],y[61]);
and and2942(ip_45_62,x[45],y[62]);
and and2943(ip_45_63,x[45],y[63]);
and and2944(ip_46_0,x[46],y[0]);
and and2945(ip_46_1,x[46],y[1]);
and and2946(ip_46_2,x[46],y[2]);
and and2947(ip_46_3,x[46],y[3]);
and and2948(ip_46_4,x[46],y[4]);
and and2949(ip_46_5,x[46],y[5]);
and and2950(ip_46_6,x[46],y[6]);
and and2951(ip_46_7,x[46],y[7]);
and and2952(ip_46_8,x[46],y[8]);
and and2953(ip_46_9,x[46],y[9]);
and and2954(ip_46_10,x[46],y[10]);
and and2955(ip_46_11,x[46],y[11]);
and and2956(ip_46_12,x[46],y[12]);
and and2957(ip_46_13,x[46],y[13]);
and and2958(ip_46_14,x[46],y[14]);
and and2959(ip_46_15,x[46],y[15]);
and and2960(ip_46_16,x[46],y[16]);
and and2961(ip_46_17,x[46],y[17]);
and and2962(ip_46_18,x[46],y[18]);
and and2963(ip_46_19,x[46],y[19]);
and and2964(ip_46_20,x[46],y[20]);
and and2965(ip_46_21,x[46],y[21]);
and and2966(ip_46_22,x[46],y[22]);
and and2967(ip_46_23,x[46],y[23]);
and and2968(ip_46_24,x[46],y[24]);
and and2969(ip_46_25,x[46],y[25]);
and and2970(ip_46_26,x[46],y[26]);
and and2971(ip_46_27,x[46],y[27]);
and and2972(ip_46_28,x[46],y[28]);
and and2973(ip_46_29,x[46],y[29]);
and and2974(ip_46_30,x[46],y[30]);
and and2975(ip_46_31,x[46],y[31]);
and and2976(ip_46_32,x[46],y[32]);
and and2977(ip_46_33,x[46],y[33]);
and and2978(ip_46_34,x[46],y[34]);
and and2979(ip_46_35,x[46],y[35]);
and and2980(ip_46_36,x[46],y[36]);
and and2981(ip_46_37,x[46],y[37]);
and and2982(ip_46_38,x[46],y[38]);
and and2983(ip_46_39,x[46],y[39]);
and and2984(ip_46_40,x[46],y[40]);
and and2985(ip_46_41,x[46],y[41]);
and and2986(ip_46_42,x[46],y[42]);
and and2987(ip_46_43,x[46],y[43]);
and and2988(ip_46_44,x[46],y[44]);
and and2989(ip_46_45,x[46],y[45]);
and and2990(ip_46_46,x[46],y[46]);
and and2991(ip_46_47,x[46],y[47]);
and and2992(ip_46_48,x[46],y[48]);
and and2993(ip_46_49,x[46],y[49]);
and and2994(ip_46_50,x[46],y[50]);
and and2995(ip_46_51,x[46],y[51]);
and and2996(ip_46_52,x[46],y[52]);
and and2997(ip_46_53,x[46],y[53]);
and and2998(ip_46_54,x[46],y[54]);
and and2999(ip_46_55,x[46],y[55]);
and and3000(ip_46_56,x[46],y[56]);
and and3001(ip_46_57,x[46],y[57]);
and and3002(ip_46_58,x[46],y[58]);
and and3003(ip_46_59,x[46],y[59]);
and and3004(ip_46_60,x[46],y[60]);
and and3005(ip_46_61,x[46],y[61]);
and and3006(ip_46_62,x[46],y[62]);
and and3007(ip_46_63,x[46],y[63]);
and and3008(ip_47_0,x[47],y[0]);
and and3009(ip_47_1,x[47],y[1]);
and and3010(ip_47_2,x[47],y[2]);
and and3011(ip_47_3,x[47],y[3]);
and and3012(ip_47_4,x[47],y[4]);
and and3013(ip_47_5,x[47],y[5]);
and and3014(ip_47_6,x[47],y[6]);
and and3015(ip_47_7,x[47],y[7]);
and and3016(ip_47_8,x[47],y[8]);
and and3017(ip_47_9,x[47],y[9]);
and and3018(ip_47_10,x[47],y[10]);
and and3019(ip_47_11,x[47],y[11]);
and and3020(ip_47_12,x[47],y[12]);
and and3021(ip_47_13,x[47],y[13]);
and and3022(ip_47_14,x[47],y[14]);
and and3023(ip_47_15,x[47],y[15]);
and and3024(ip_47_16,x[47],y[16]);
and and3025(ip_47_17,x[47],y[17]);
and and3026(ip_47_18,x[47],y[18]);
and and3027(ip_47_19,x[47],y[19]);
and and3028(ip_47_20,x[47],y[20]);
and and3029(ip_47_21,x[47],y[21]);
and and3030(ip_47_22,x[47],y[22]);
and and3031(ip_47_23,x[47],y[23]);
and and3032(ip_47_24,x[47],y[24]);
and and3033(ip_47_25,x[47],y[25]);
and and3034(ip_47_26,x[47],y[26]);
and and3035(ip_47_27,x[47],y[27]);
and and3036(ip_47_28,x[47],y[28]);
and and3037(ip_47_29,x[47],y[29]);
and and3038(ip_47_30,x[47],y[30]);
and and3039(ip_47_31,x[47],y[31]);
and and3040(ip_47_32,x[47],y[32]);
and and3041(ip_47_33,x[47],y[33]);
and and3042(ip_47_34,x[47],y[34]);
and and3043(ip_47_35,x[47],y[35]);
and and3044(ip_47_36,x[47],y[36]);
and and3045(ip_47_37,x[47],y[37]);
and and3046(ip_47_38,x[47],y[38]);
and and3047(ip_47_39,x[47],y[39]);
and and3048(ip_47_40,x[47],y[40]);
and and3049(ip_47_41,x[47],y[41]);
and and3050(ip_47_42,x[47],y[42]);
and and3051(ip_47_43,x[47],y[43]);
and and3052(ip_47_44,x[47],y[44]);
and and3053(ip_47_45,x[47],y[45]);
and and3054(ip_47_46,x[47],y[46]);
and and3055(ip_47_47,x[47],y[47]);
and and3056(ip_47_48,x[47],y[48]);
and and3057(ip_47_49,x[47],y[49]);
and and3058(ip_47_50,x[47],y[50]);
and and3059(ip_47_51,x[47],y[51]);
and and3060(ip_47_52,x[47],y[52]);
and and3061(ip_47_53,x[47],y[53]);
and and3062(ip_47_54,x[47],y[54]);
and and3063(ip_47_55,x[47],y[55]);
and and3064(ip_47_56,x[47],y[56]);
and and3065(ip_47_57,x[47],y[57]);
and and3066(ip_47_58,x[47],y[58]);
and and3067(ip_47_59,x[47],y[59]);
and and3068(ip_47_60,x[47],y[60]);
and and3069(ip_47_61,x[47],y[61]);
and and3070(ip_47_62,x[47],y[62]);
and and3071(ip_47_63,x[47],y[63]);
and and3072(ip_48_0,x[48],y[0]);
and and3073(ip_48_1,x[48],y[1]);
and and3074(ip_48_2,x[48],y[2]);
and and3075(ip_48_3,x[48],y[3]);
and and3076(ip_48_4,x[48],y[4]);
and and3077(ip_48_5,x[48],y[5]);
and and3078(ip_48_6,x[48],y[6]);
and and3079(ip_48_7,x[48],y[7]);
and and3080(ip_48_8,x[48],y[8]);
and and3081(ip_48_9,x[48],y[9]);
and and3082(ip_48_10,x[48],y[10]);
and and3083(ip_48_11,x[48],y[11]);
and and3084(ip_48_12,x[48],y[12]);
and and3085(ip_48_13,x[48],y[13]);
and and3086(ip_48_14,x[48],y[14]);
and and3087(ip_48_15,x[48],y[15]);
and and3088(ip_48_16,x[48],y[16]);
and and3089(ip_48_17,x[48],y[17]);
and and3090(ip_48_18,x[48],y[18]);
and and3091(ip_48_19,x[48],y[19]);
and and3092(ip_48_20,x[48],y[20]);
and and3093(ip_48_21,x[48],y[21]);
and and3094(ip_48_22,x[48],y[22]);
and and3095(ip_48_23,x[48],y[23]);
and and3096(ip_48_24,x[48],y[24]);
and and3097(ip_48_25,x[48],y[25]);
and and3098(ip_48_26,x[48],y[26]);
and and3099(ip_48_27,x[48],y[27]);
and and3100(ip_48_28,x[48],y[28]);
and and3101(ip_48_29,x[48],y[29]);
and and3102(ip_48_30,x[48],y[30]);
and and3103(ip_48_31,x[48],y[31]);
and and3104(ip_48_32,x[48],y[32]);
and and3105(ip_48_33,x[48],y[33]);
and and3106(ip_48_34,x[48],y[34]);
and and3107(ip_48_35,x[48],y[35]);
and and3108(ip_48_36,x[48],y[36]);
and and3109(ip_48_37,x[48],y[37]);
and and3110(ip_48_38,x[48],y[38]);
and and3111(ip_48_39,x[48],y[39]);
and and3112(ip_48_40,x[48],y[40]);
and and3113(ip_48_41,x[48],y[41]);
and and3114(ip_48_42,x[48],y[42]);
and and3115(ip_48_43,x[48],y[43]);
and and3116(ip_48_44,x[48],y[44]);
and and3117(ip_48_45,x[48],y[45]);
and and3118(ip_48_46,x[48],y[46]);
and and3119(ip_48_47,x[48],y[47]);
and and3120(ip_48_48,x[48],y[48]);
and and3121(ip_48_49,x[48],y[49]);
and and3122(ip_48_50,x[48],y[50]);
and and3123(ip_48_51,x[48],y[51]);
and and3124(ip_48_52,x[48],y[52]);
and and3125(ip_48_53,x[48],y[53]);
and and3126(ip_48_54,x[48],y[54]);
and and3127(ip_48_55,x[48],y[55]);
and and3128(ip_48_56,x[48],y[56]);
and and3129(ip_48_57,x[48],y[57]);
and and3130(ip_48_58,x[48],y[58]);
and and3131(ip_48_59,x[48],y[59]);
and and3132(ip_48_60,x[48],y[60]);
and and3133(ip_48_61,x[48],y[61]);
and and3134(ip_48_62,x[48],y[62]);
and and3135(ip_48_63,x[48],y[63]);
and and3136(ip_49_0,x[49],y[0]);
and and3137(ip_49_1,x[49],y[1]);
and and3138(ip_49_2,x[49],y[2]);
and and3139(ip_49_3,x[49],y[3]);
and and3140(ip_49_4,x[49],y[4]);
and and3141(ip_49_5,x[49],y[5]);
and and3142(ip_49_6,x[49],y[6]);
and and3143(ip_49_7,x[49],y[7]);
and and3144(ip_49_8,x[49],y[8]);
and and3145(ip_49_9,x[49],y[9]);
and and3146(ip_49_10,x[49],y[10]);
and and3147(ip_49_11,x[49],y[11]);
and and3148(ip_49_12,x[49],y[12]);
and and3149(ip_49_13,x[49],y[13]);
and and3150(ip_49_14,x[49],y[14]);
and and3151(ip_49_15,x[49],y[15]);
and and3152(ip_49_16,x[49],y[16]);
and and3153(ip_49_17,x[49],y[17]);
and and3154(ip_49_18,x[49],y[18]);
and and3155(ip_49_19,x[49],y[19]);
and and3156(ip_49_20,x[49],y[20]);
and and3157(ip_49_21,x[49],y[21]);
and and3158(ip_49_22,x[49],y[22]);
and and3159(ip_49_23,x[49],y[23]);
and and3160(ip_49_24,x[49],y[24]);
and and3161(ip_49_25,x[49],y[25]);
and and3162(ip_49_26,x[49],y[26]);
and and3163(ip_49_27,x[49],y[27]);
and and3164(ip_49_28,x[49],y[28]);
and and3165(ip_49_29,x[49],y[29]);
and and3166(ip_49_30,x[49],y[30]);
and and3167(ip_49_31,x[49],y[31]);
and and3168(ip_49_32,x[49],y[32]);
and and3169(ip_49_33,x[49],y[33]);
and and3170(ip_49_34,x[49],y[34]);
and and3171(ip_49_35,x[49],y[35]);
and and3172(ip_49_36,x[49],y[36]);
and and3173(ip_49_37,x[49],y[37]);
and and3174(ip_49_38,x[49],y[38]);
and and3175(ip_49_39,x[49],y[39]);
and and3176(ip_49_40,x[49],y[40]);
and and3177(ip_49_41,x[49],y[41]);
and and3178(ip_49_42,x[49],y[42]);
and and3179(ip_49_43,x[49],y[43]);
and and3180(ip_49_44,x[49],y[44]);
and and3181(ip_49_45,x[49],y[45]);
and and3182(ip_49_46,x[49],y[46]);
and and3183(ip_49_47,x[49],y[47]);
and and3184(ip_49_48,x[49],y[48]);
and and3185(ip_49_49,x[49],y[49]);
and and3186(ip_49_50,x[49],y[50]);
and and3187(ip_49_51,x[49],y[51]);
and and3188(ip_49_52,x[49],y[52]);
and and3189(ip_49_53,x[49],y[53]);
and and3190(ip_49_54,x[49],y[54]);
and and3191(ip_49_55,x[49],y[55]);
and and3192(ip_49_56,x[49],y[56]);
and and3193(ip_49_57,x[49],y[57]);
and and3194(ip_49_58,x[49],y[58]);
and and3195(ip_49_59,x[49],y[59]);
and and3196(ip_49_60,x[49],y[60]);
and and3197(ip_49_61,x[49],y[61]);
and and3198(ip_49_62,x[49],y[62]);
and and3199(ip_49_63,x[49],y[63]);
and and3200(ip_50_0,x[50],y[0]);
and and3201(ip_50_1,x[50],y[1]);
and and3202(ip_50_2,x[50],y[2]);
and and3203(ip_50_3,x[50],y[3]);
and and3204(ip_50_4,x[50],y[4]);
and and3205(ip_50_5,x[50],y[5]);
and and3206(ip_50_6,x[50],y[6]);
and and3207(ip_50_7,x[50],y[7]);
and and3208(ip_50_8,x[50],y[8]);
and and3209(ip_50_9,x[50],y[9]);
and and3210(ip_50_10,x[50],y[10]);
and and3211(ip_50_11,x[50],y[11]);
and and3212(ip_50_12,x[50],y[12]);
and and3213(ip_50_13,x[50],y[13]);
and and3214(ip_50_14,x[50],y[14]);
and and3215(ip_50_15,x[50],y[15]);
and and3216(ip_50_16,x[50],y[16]);
and and3217(ip_50_17,x[50],y[17]);
and and3218(ip_50_18,x[50],y[18]);
and and3219(ip_50_19,x[50],y[19]);
and and3220(ip_50_20,x[50],y[20]);
and and3221(ip_50_21,x[50],y[21]);
and and3222(ip_50_22,x[50],y[22]);
and and3223(ip_50_23,x[50],y[23]);
and and3224(ip_50_24,x[50],y[24]);
and and3225(ip_50_25,x[50],y[25]);
and and3226(ip_50_26,x[50],y[26]);
and and3227(ip_50_27,x[50],y[27]);
and and3228(ip_50_28,x[50],y[28]);
and and3229(ip_50_29,x[50],y[29]);
and and3230(ip_50_30,x[50],y[30]);
and and3231(ip_50_31,x[50],y[31]);
and and3232(ip_50_32,x[50],y[32]);
and and3233(ip_50_33,x[50],y[33]);
and and3234(ip_50_34,x[50],y[34]);
and and3235(ip_50_35,x[50],y[35]);
and and3236(ip_50_36,x[50],y[36]);
and and3237(ip_50_37,x[50],y[37]);
and and3238(ip_50_38,x[50],y[38]);
and and3239(ip_50_39,x[50],y[39]);
and and3240(ip_50_40,x[50],y[40]);
and and3241(ip_50_41,x[50],y[41]);
and and3242(ip_50_42,x[50],y[42]);
and and3243(ip_50_43,x[50],y[43]);
and and3244(ip_50_44,x[50],y[44]);
and and3245(ip_50_45,x[50],y[45]);
and and3246(ip_50_46,x[50],y[46]);
and and3247(ip_50_47,x[50],y[47]);
and and3248(ip_50_48,x[50],y[48]);
and and3249(ip_50_49,x[50],y[49]);
and and3250(ip_50_50,x[50],y[50]);
and and3251(ip_50_51,x[50],y[51]);
and and3252(ip_50_52,x[50],y[52]);
and and3253(ip_50_53,x[50],y[53]);
and and3254(ip_50_54,x[50],y[54]);
and and3255(ip_50_55,x[50],y[55]);
and and3256(ip_50_56,x[50],y[56]);
and and3257(ip_50_57,x[50],y[57]);
and and3258(ip_50_58,x[50],y[58]);
and and3259(ip_50_59,x[50],y[59]);
and and3260(ip_50_60,x[50],y[60]);
and and3261(ip_50_61,x[50],y[61]);
and and3262(ip_50_62,x[50],y[62]);
and and3263(ip_50_63,x[50],y[63]);
and and3264(ip_51_0,x[51],y[0]);
and and3265(ip_51_1,x[51],y[1]);
and and3266(ip_51_2,x[51],y[2]);
and and3267(ip_51_3,x[51],y[3]);
and and3268(ip_51_4,x[51],y[4]);
and and3269(ip_51_5,x[51],y[5]);
and and3270(ip_51_6,x[51],y[6]);
and and3271(ip_51_7,x[51],y[7]);
and and3272(ip_51_8,x[51],y[8]);
and and3273(ip_51_9,x[51],y[9]);
and and3274(ip_51_10,x[51],y[10]);
and and3275(ip_51_11,x[51],y[11]);
and and3276(ip_51_12,x[51],y[12]);
and and3277(ip_51_13,x[51],y[13]);
and and3278(ip_51_14,x[51],y[14]);
and and3279(ip_51_15,x[51],y[15]);
and and3280(ip_51_16,x[51],y[16]);
and and3281(ip_51_17,x[51],y[17]);
and and3282(ip_51_18,x[51],y[18]);
and and3283(ip_51_19,x[51],y[19]);
and and3284(ip_51_20,x[51],y[20]);
and and3285(ip_51_21,x[51],y[21]);
and and3286(ip_51_22,x[51],y[22]);
and and3287(ip_51_23,x[51],y[23]);
and and3288(ip_51_24,x[51],y[24]);
and and3289(ip_51_25,x[51],y[25]);
and and3290(ip_51_26,x[51],y[26]);
and and3291(ip_51_27,x[51],y[27]);
and and3292(ip_51_28,x[51],y[28]);
and and3293(ip_51_29,x[51],y[29]);
and and3294(ip_51_30,x[51],y[30]);
and and3295(ip_51_31,x[51],y[31]);
and and3296(ip_51_32,x[51],y[32]);
and and3297(ip_51_33,x[51],y[33]);
and and3298(ip_51_34,x[51],y[34]);
and and3299(ip_51_35,x[51],y[35]);
and and3300(ip_51_36,x[51],y[36]);
and and3301(ip_51_37,x[51],y[37]);
and and3302(ip_51_38,x[51],y[38]);
and and3303(ip_51_39,x[51],y[39]);
and and3304(ip_51_40,x[51],y[40]);
and and3305(ip_51_41,x[51],y[41]);
and and3306(ip_51_42,x[51],y[42]);
and and3307(ip_51_43,x[51],y[43]);
and and3308(ip_51_44,x[51],y[44]);
and and3309(ip_51_45,x[51],y[45]);
and and3310(ip_51_46,x[51],y[46]);
and and3311(ip_51_47,x[51],y[47]);
and and3312(ip_51_48,x[51],y[48]);
and and3313(ip_51_49,x[51],y[49]);
and and3314(ip_51_50,x[51],y[50]);
and and3315(ip_51_51,x[51],y[51]);
and and3316(ip_51_52,x[51],y[52]);
and and3317(ip_51_53,x[51],y[53]);
and and3318(ip_51_54,x[51],y[54]);
and and3319(ip_51_55,x[51],y[55]);
and and3320(ip_51_56,x[51],y[56]);
and and3321(ip_51_57,x[51],y[57]);
and and3322(ip_51_58,x[51],y[58]);
and and3323(ip_51_59,x[51],y[59]);
and and3324(ip_51_60,x[51],y[60]);
and and3325(ip_51_61,x[51],y[61]);
and and3326(ip_51_62,x[51],y[62]);
and and3327(ip_51_63,x[51],y[63]);
and and3328(ip_52_0,x[52],y[0]);
and and3329(ip_52_1,x[52],y[1]);
and and3330(ip_52_2,x[52],y[2]);
and and3331(ip_52_3,x[52],y[3]);
and and3332(ip_52_4,x[52],y[4]);
and and3333(ip_52_5,x[52],y[5]);
and and3334(ip_52_6,x[52],y[6]);
and and3335(ip_52_7,x[52],y[7]);
and and3336(ip_52_8,x[52],y[8]);
and and3337(ip_52_9,x[52],y[9]);
and and3338(ip_52_10,x[52],y[10]);
and and3339(ip_52_11,x[52],y[11]);
and and3340(ip_52_12,x[52],y[12]);
and and3341(ip_52_13,x[52],y[13]);
and and3342(ip_52_14,x[52],y[14]);
and and3343(ip_52_15,x[52],y[15]);
and and3344(ip_52_16,x[52],y[16]);
and and3345(ip_52_17,x[52],y[17]);
and and3346(ip_52_18,x[52],y[18]);
and and3347(ip_52_19,x[52],y[19]);
and and3348(ip_52_20,x[52],y[20]);
and and3349(ip_52_21,x[52],y[21]);
and and3350(ip_52_22,x[52],y[22]);
and and3351(ip_52_23,x[52],y[23]);
and and3352(ip_52_24,x[52],y[24]);
and and3353(ip_52_25,x[52],y[25]);
and and3354(ip_52_26,x[52],y[26]);
and and3355(ip_52_27,x[52],y[27]);
and and3356(ip_52_28,x[52],y[28]);
and and3357(ip_52_29,x[52],y[29]);
and and3358(ip_52_30,x[52],y[30]);
and and3359(ip_52_31,x[52],y[31]);
and and3360(ip_52_32,x[52],y[32]);
and and3361(ip_52_33,x[52],y[33]);
and and3362(ip_52_34,x[52],y[34]);
and and3363(ip_52_35,x[52],y[35]);
and and3364(ip_52_36,x[52],y[36]);
and and3365(ip_52_37,x[52],y[37]);
and and3366(ip_52_38,x[52],y[38]);
and and3367(ip_52_39,x[52],y[39]);
and and3368(ip_52_40,x[52],y[40]);
and and3369(ip_52_41,x[52],y[41]);
and and3370(ip_52_42,x[52],y[42]);
and and3371(ip_52_43,x[52],y[43]);
and and3372(ip_52_44,x[52],y[44]);
and and3373(ip_52_45,x[52],y[45]);
and and3374(ip_52_46,x[52],y[46]);
and and3375(ip_52_47,x[52],y[47]);
and and3376(ip_52_48,x[52],y[48]);
and and3377(ip_52_49,x[52],y[49]);
and and3378(ip_52_50,x[52],y[50]);
and and3379(ip_52_51,x[52],y[51]);
and and3380(ip_52_52,x[52],y[52]);
and and3381(ip_52_53,x[52],y[53]);
and and3382(ip_52_54,x[52],y[54]);
and and3383(ip_52_55,x[52],y[55]);
and and3384(ip_52_56,x[52],y[56]);
and and3385(ip_52_57,x[52],y[57]);
and and3386(ip_52_58,x[52],y[58]);
and and3387(ip_52_59,x[52],y[59]);
and and3388(ip_52_60,x[52],y[60]);
and and3389(ip_52_61,x[52],y[61]);
and and3390(ip_52_62,x[52],y[62]);
and and3391(ip_52_63,x[52],y[63]);
and and3392(ip_53_0,x[53],y[0]);
and and3393(ip_53_1,x[53],y[1]);
and and3394(ip_53_2,x[53],y[2]);
and and3395(ip_53_3,x[53],y[3]);
and and3396(ip_53_4,x[53],y[4]);
and and3397(ip_53_5,x[53],y[5]);
and and3398(ip_53_6,x[53],y[6]);
and and3399(ip_53_7,x[53],y[7]);
and and3400(ip_53_8,x[53],y[8]);
and and3401(ip_53_9,x[53],y[9]);
and and3402(ip_53_10,x[53],y[10]);
and and3403(ip_53_11,x[53],y[11]);
and and3404(ip_53_12,x[53],y[12]);
and and3405(ip_53_13,x[53],y[13]);
and and3406(ip_53_14,x[53],y[14]);
and and3407(ip_53_15,x[53],y[15]);
and and3408(ip_53_16,x[53],y[16]);
and and3409(ip_53_17,x[53],y[17]);
and and3410(ip_53_18,x[53],y[18]);
and and3411(ip_53_19,x[53],y[19]);
and and3412(ip_53_20,x[53],y[20]);
and and3413(ip_53_21,x[53],y[21]);
and and3414(ip_53_22,x[53],y[22]);
and and3415(ip_53_23,x[53],y[23]);
and and3416(ip_53_24,x[53],y[24]);
and and3417(ip_53_25,x[53],y[25]);
and and3418(ip_53_26,x[53],y[26]);
and and3419(ip_53_27,x[53],y[27]);
and and3420(ip_53_28,x[53],y[28]);
and and3421(ip_53_29,x[53],y[29]);
and and3422(ip_53_30,x[53],y[30]);
and and3423(ip_53_31,x[53],y[31]);
and and3424(ip_53_32,x[53],y[32]);
and and3425(ip_53_33,x[53],y[33]);
and and3426(ip_53_34,x[53],y[34]);
and and3427(ip_53_35,x[53],y[35]);
and and3428(ip_53_36,x[53],y[36]);
and and3429(ip_53_37,x[53],y[37]);
and and3430(ip_53_38,x[53],y[38]);
and and3431(ip_53_39,x[53],y[39]);
and and3432(ip_53_40,x[53],y[40]);
and and3433(ip_53_41,x[53],y[41]);
and and3434(ip_53_42,x[53],y[42]);
and and3435(ip_53_43,x[53],y[43]);
and and3436(ip_53_44,x[53],y[44]);
and and3437(ip_53_45,x[53],y[45]);
and and3438(ip_53_46,x[53],y[46]);
and and3439(ip_53_47,x[53],y[47]);
and and3440(ip_53_48,x[53],y[48]);
and and3441(ip_53_49,x[53],y[49]);
and and3442(ip_53_50,x[53],y[50]);
and and3443(ip_53_51,x[53],y[51]);
and and3444(ip_53_52,x[53],y[52]);
and and3445(ip_53_53,x[53],y[53]);
and and3446(ip_53_54,x[53],y[54]);
and and3447(ip_53_55,x[53],y[55]);
and and3448(ip_53_56,x[53],y[56]);
and and3449(ip_53_57,x[53],y[57]);
and and3450(ip_53_58,x[53],y[58]);
and and3451(ip_53_59,x[53],y[59]);
and and3452(ip_53_60,x[53],y[60]);
and and3453(ip_53_61,x[53],y[61]);
and and3454(ip_53_62,x[53],y[62]);
and and3455(ip_53_63,x[53],y[63]);
and and3456(ip_54_0,x[54],y[0]);
and and3457(ip_54_1,x[54],y[1]);
and and3458(ip_54_2,x[54],y[2]);
and and3459(ip_54_3,x[54],y[3]);
and and3460(ip_54_4,x[54],y[4]);
and and3461(ip_54_5,x[54],y[5]);
and and3462(ip_54_6,x[54],y[6]);
and and3463(ip_54_7,x[54],y[7]);
and and3464(ip_54_8,x[54],y[8]);
and and3465(ip_54_9,x[54],y[9]);
and and3466(ip_54_10,x[54],y[10]);
and and3467(ip_54_11,x[54],y[11]);
and and3468(ip_54_12,x[54],y[12]);
and and3469(ip_54_13,x[54],y[13]);
and and3470(ip_54_14,x[54],y[14]);
and and3471(ip_54_15,x[54],y[15]);
and and3472(ip_54_16,x[54],y[16]);
and and3473(ip_54_17,x[54],y[17]);
and and3474(ip_54_18,x[54],y[18]);
and and3475(ip_54_19,x[54],y[19]);
and and3476(ip_54_20,x[54],y[20]);
and and3477(ip_54_21,x[54],y[21]);
and and3478(ip_54_22,x[54],y[22]);
and and3479(ip_54_23,x[54],y[23]);
and and3480(ip_54_24,x[54],y[24]);
and and3481(ip_54_25,x[54],y[25]);
and and3482(ip_54_26,x[54],y[26]);
and and3483(ip_54_27,x[54],y[27]);
and and3484(ip_54_28,x[54],y[28]);
and and3485(ip_54_29,x[54],y[29]);
and and3486(ip_54_30,x[54],y[30]);
and and3487(ip_54_31,x[54],y[31]);
and and3488(ip_54_32,x[54],y[32]);
and and3489(ip_54_33,x[54],y[33]);
and and3490(ip_54_34,x[54],y[34]);
and and3491(ip_54_35,x[54],y[35]);
and and3492(ip_54_36,x[54],y[36]);
and and3493(ip_54_37,x[54],y[37]);
and and3494(ip_54_38,x[54],y[38]);
and and3495(ip_54_39,x[54],y[39]);
and and3496(ip_54_40,x[54],y[40]);
and and3497(ip_54_41,x[54],y[41]);
and and3498(ip_54_42,x[54],y[42]);
and and3499(ip_54_43,x[54],y[43]);
and and3500(ip_54_44,x[54],y[44]);
and and3501(ip_54_45,x[54],y[45]);
and and3502(ip_54_46,x[54],y[46]);
and and3503(ip_54_47,x[54],y[47]);
and and3504(ip_54_48,x[54],y[48]);
and and3505(ip_54_49,x[54],y[49]);
and and3506(ip_54_50,x[54],y[50]);
and and3507(ip_54_51,x[54],y[51]);
and and3508(ip_54_52,x[54],y[52]);
and and3509(ip_54_53,x[54],y[53]);
and and3510(ip_54_54,x[54],y[54]);
and and3511(ip_54_55,x[54],y[55]);
and and3512(ip_54_56,x[54],y[56]);
and and3513(ip_54_57,x[54],y[57]);
and and3514(ip_54_58,x[54],y[58]);
and and3515(ip_54_59,x[54],y[59]);
and and3516(ip_54_60,x[54],y[60]);
and and3517(ip_54_61,x[54],y[61]);
and and3518(ip_54_62,x[54],y[62]);
and and3519(ip_54_63,x[54],y[63]);
and and3520(ip_55_0,x[55],y[0]);
and and3521(ip_55_1,x[55],y[1]);
and and3522(ip_55_2,x[55],y[2]);
and and3523(ip_55_3,x[55],y[3]);
and and3524(ip_55_4,x[55],y[4]);
and and3525(ip_55_5,x[55],y[5]);
and and3526(ip_55_6,x[55],y[6]);
and and3527(ip_55_7,x[55],y[7]);
and and3528(ip_55_8,x[55],y[8]);
and and3529(ip_55_9,x[55],y[9]);
and and3530(ip_55_10,x[55],y[10]);
and and3531(ip_55_11,x[55],y[11]);
and and3532(ip_55_12,x[55],y[12]);
and and3533(ip_55_13,x[55],y[13]);
and and3534(ip_55_14,x[55],y[14]);
and and3535(ip_55_15,x[55],y[15]);
and and3536(ip_55_16,x[55],y[16]);
and and3537(ip_55_17,x[55],y[17]);
and and3538(ip_55_18,x[55],y[18]);
and and3539(ip_55_19,x[55],y[19]);
and and3540(ip_55_20,x[55],y[20]);
and and3541(ip_55_21,x[55],y[21]);
and and3542(ip_55_22,x[55],y[22]);
and and3543(ip_55_23,x[55],y[23]);
and and3544(ip_55_24,x[55],y[24]);
and and3545(ip_55_25,x[55],y[25]);
and and3546(ip_55_26,x[55],y[26]);
and and3547(ip_55_27,x[55],y[27]);
and and3548(ip_55_28,x[55],y[28]);
and and3549(ip_55_29,x[55],y[29]);
and and3550(ip_55_30,x[55],y[30]);
and and3551(ip_55_31,x[55],y[31]);
and and3552(ip_55_32,x[55],y[32]);
and and3553(ip_55_33,x[55],y[33]);
and and3554(ip_55_34,x[55],y[34]);
and and3555(ip_55_35,x[55],y[35]);
and and3556(ip_55_36,x[55],y[36]);
and and3557(ip_55_37,x[55],y[37]);
and and3558(ip_55_38,x[55],y[38]);
and and3559(ip_55_39,x[55],y[39]);
and and3560(ip_55_40,x[55],y[40]);
and and3561(ip_55_41,x[55],y[41]);
and and3562(ip_55_42,x[55],y[42]);
and and3563(ip_55_43,x[55],y[43]);
and and3564(ip_55_44,x[55],y[44]);
and and3565(ip_55_45,x[55],y[45]);
and and3566(ip_55_46,x[55],y[46]);
and and3567(ip_55_47,x[55],y[47]);
and and3568(ip_55_48,x[55],y[48]);
and and3569(ip_55_49,x[55],y[49]);
and and3570(ip_55_50,x[55],y[50]);
and and3571(ip_55_51,x[55],y[51]);
and and3572(ip_55_52,x[55],y[52]);
and and3573(ip_55_53,x[55],y[53]);
and and3574(ip_55_54,x[55],y[54]);
and and3575(ip_55_55,x[55],y[55]);
and and3576(ip_55_56,x[55],y[56]);
and and3577(ip_55_57,x[55],y[57]);
and and3578(ip_55_58,x[55],y[58]);
and and3579(ip_55_59,x[55],y[59]);
and and3580(ip_55_60,x[55],y[60]);
and and3581(ip_55_61,x[55],y[61]);
and and3582(ip_55_62,x[55],y[62]);
and and3583(ip_55_63,x[55],y[63]);
and and3584(ip_56_0,x[56],y[0]);
and and3585(ip_56_1,x[56],y[1]);
and and3586(ip_56_2,x[56],y[2]);
and and3587(ip_56_3,x[56],y[3]);
and and3588(ip_56_4,x[56],y[4]);
and and3589(ip_56_5,x[56],y[5]);
and and3590(ip_56_6,x[56],y[6]);
and and3591(ip_56_7,x[56],y[7]);
and and3592(ip_56_8,x[56],y[8]);
and and3593(ip_56_9,x[56],y[9]);
and and3594(ip_56_10,x[56],y[10]);
and and3595(ip_56_11,x[56],y[11]);
and and3596(ip_56_12,x[56],y[12]);
and and3597(ip_56_13,x[56],y[13]);
and and3598(ip_56_14,x[56],y[14]);
and and3599(ip_56_15,x[56],y[15]);
and and3600(ip_56_16,x[56],y[16]);
and and3601(ip_56_17,x[56],y[17]);
and and3602(ip_56_18,x[56],y[18]);
and and3603(ip_56_19,x[56],y[19]);
and and3604(ip_56_20,x[56],y[20]);
and and3605(ip_56_21,x[56],y[21]);
and and3606(ip_56_22,x[56],y[22]);
and and3607(ip_56_23,x[56],y[23]);
and and3608(ip_56_24,x[56],y[24]);
and and3609(ip_56_25,x[56],y[25]);
and and3610(ip_56_26,x[56],y[26]);
and and3611(ip_56_27,x[56],y[27]);
and and3612(ip_56_28,x[56],y[28]);
and and3613(ip_56_29,x[56],y[29]);
and and3614(ip_56_30,x[56],y[30]);
and and3615(ip_56_31,x[56],y[31]);
and and3616(ip_56_32,x[56],y[32]);
and and3617(ip_56_33,x[56],y[33]);
and and3618(ip_56_34,x[56],y[34]);
and and3619(ip_56_35,x[56],y[35]);
and and3620(ip_56_36,x[56],y[36]);
and and3621(ip_56_37,x[56],y[37]);
and and3622(ip_56_38,x[56],y[38]);
and and3623(ip_56_39,x[56],y[39]);
and and3624(ip_56_40,x[56],y[40]);
and and3625(ip_56_41,x[56],y[41]);
and and3626(ip_56_42,x[56],y[42]);
and and3627(ip_56_43,x[56],y[43]);
and and3628(ip_56_44,x[56],y[44]);
and and3629(ip_56_45,x[56],y[45]);
and and3630(ip_56_46,x[56],y[46]);
and and3631(ip_56_47,x[56],y[47]);
and and3632(ip_56_48,x[56],y[48]);
and and3633(ip_56_49,x[56],y[49]);
and and3634(ip_56_50,x[56],y[50]);
and and3635(ip_56_51,x[56],y[51]);
and and3636(ip_56_52,x[56],y[52]);
and and3637(ip_56_53,x[56],y[53]);
and and3638(ip_56_54,x[56],y[54]);
and and3639(ip_56_55,x[56],y[55]);
and and3640(ip_56_56,x[56],y[56]);
and and3641(ip_56_57,x[56],y[57]);
and and3642(ip_56_58,x[56],y[58]);
and and3643(ip_56_59,x[56],y[59]);
and and3644(ip_56_60,x[56],y[60]);
and and3645(ip_56_61,x[56],y[61]);
and and3646(ip_56_62,x[56],y[62]);
and and3647(ip_56_63,x[56],y[63]);
and and3648(ip_57_0,x[57],y[0]);
and and3649(ip_57_1,x[57],y[1]);
and and3650(ip_57_2,x[57],y[2]);
and and3651(ip_57_3,x[57],y[3]);
and and3652(ip_57_4,x[57],y[4]);
and and3653(ip_57_5,x[57],y[5]);
and and3654(ip_57_6,x[57],y[6]);
and and3655(ip_57_7,x[57],y[7]);
and and3656(ip_57_8,x[57],y[8]);
and and3657(ip_57_9,x[57],y[9]);
and and3658(ip_57_10,x[57],y[10]);
and and3659(ip_57_11,x[57],y[11]);
and and3660(ip_57_12,x[57],y[12]);
and and3661(ip_57_13,x[57],y[13]);
and and3662(ip_57_14,x[57],y[14]);
and and3663(ip_57_15,x[57],y[15]);
and and3664(ip_57_16,x[57],y[16]);
and and3665(ip_57_17,x[57],y[17]);
and and3666(ip_57_18,x[57],y[18]);
and and3667(ip_57_19,x[57],y[19]);
and and3668(ip_57_20,x[57],y[20]);
and and3669(ip_57_21,x[57],y[21]);
and and3670(ip_57_22,x[57],y[22]);
and and3671(ip_57_23,x[57],y[23]);
and and3672(ip_57_24,x[57],y[24]);
and and3673(ip_57_25,x[57],y[25]);
and and3674(ip_57_26,x[57],y[26]);
and and3675(ip_57_27,x[57],y[27]);
and and3676(ip_57_28,x[57],y[28]);
and and3677(ip_57_29,x[57],y[29]);
and and3678(ip_57_30,x[57],y[30]);
and and3679(ip_57_31,x[57],y[31]);
and and3680(ip_57_32,x[57],y[32]);
and and3681(ip_57_33,x[57],y[33]);
and and3682(ip_57_34,x[57],y[34]);
and and3683(ip_57_35,x[57],y[35]);
and and3684(ip_57_36,x[57],y[36]);
and and3685(ip_57_37,x[57],y[37]);
and and3686(ip_57_38,x[57],y[38]);
and and3687(ip_57_39,x[57],y[39]);
and and3688(ip_57_40,x[57],y[40]);
and and3689(ip_57_41,x[57],y[41]);
and and3690(ip_57_42,x[57],y[42]);
and and3691(ip_57_43,x[57],y[43]);
and and3692(ip_57_44,x[57],y[44]);
and and3693(ip_57_45,x[57],y[45]);
and and3694(ip_57_46,x[57],y[46]);
and and3695(ip_57_47,x[57],y[47]);
and and3696(ip_57_48,x[57],y[48]);
and and3697(ip_57_49,x[57],y[49]);
and and3698(ip_57_50,x[57],y[50]);
and and3699(ip_57_51,x[57],y[51]);
and and3700(ip_57_52,x[57],y[52]);
and and3701(ip_57_53,x[57],y[53]);
and and3702(ip_57_54,x[57],y[54]);
and and3703(ip_57_55,x[57],y[55]);
and and3704(ip_57_56,x[57],y[56]);
and and3705(ip_57_57,x[57],y[57]);
and and3706(ip_57_58,x[57],y[58]);
and and3707(ip_57_59,x[57],y[59]);
and and3708(ip_57_60,x[57],y[60]);
and and3709(ip_57_61,x[57],y[61]);
and and3710(ip_57_62,x[57],y[62]);
and and3711(ip_57_63,x[57],y[63]);
and and3712(ip_58_0,x[58],y[0]);
and and3713(ip_58_1,x[58],y[1]);
and and3714(ip_58_2,x[58],y[2]);
and and3715(ip_58_3,x[58],y[3]);
and and3716(ip_58_4,x[58],y[4]);
and and3717(ip_58_5,x[58],y[5]);
and and3718(ip_58_6,x[58],y[6]);
and and3719(ip_58_7,x[58],y[7]);
and and3720(ip_58_8,x[58],y[8]);
and and3721(ip_58_9,x[58],y[9]);
and and3722(ip_58_10,x[58],y[10]);
and and3723(ip_58_11,x[58],y[11]);
and and3724(ip_58_12,x[58],y[12]);
and and3725(ip_58_13,x[58],y[13]);
and and3726(ip_58_14,x[58],y[14]);
and and3727(ip_58_15,x[58],y[15]);
and and3728(ip_58_16,x[58],y[16]);
and and3729(ip_58_17,x[58],y[17]);
and and3730(ip_58_18,x[58],y[18]);
and and3731(ip_58_19,x[58],y[19]);
and and3732(ip_58_20,x[58],y[20]);
and and3733(ip_58_21,x[58],y[21]);
and and3734(ip_58_22,x[58],y[22]);
and and3735(ip_58_23,x[58],y[23]);
and and3736(ip_58_24,x[58],y[24]);
and and3737(ip_58_25,x[58],y[25]);
and and3738(ip_58_26,x[58],y[26]);
and and3739(ip_58_27,x[58],y[27]);
and and3740(ip_58_28,x[58],y[28]);
and and3741(ip_58_29,x[58],y[29]);
and and3742(ip_58_30,x[58],y[30]);
and and3743(ip_58_31,x[58],y[31]);
and and3744(ip_58_32,x[58],y[32]);
and and3745(ip_58_33,x[58],y[33]);
and and3746(ip_58_34,x[58],y[34]);
and and3747(ip_58_35,x[58],y[35]);
and and3748(ip_58_36,x[58],y[36]);
and and3749(ip_58_37,x[58],y[37]);
and and3750(ip_58_38,x[58],y[38]);
and and3751(ip_58_39,x[58],y[39]);
and and3752(ip_58_40,x[58],y[40]);
and and3753(ip_58_41,x[58],y[41]);
and and3754(ip_58_42,x[58],y[42]);
and and3755(ip_58_43,x[58],y[43]);
and and3756(ip_58_44,x[58],y[44]);
and and3757(ip_58_45,x[58],y[45]);
and and3758(ip_58_46,x[58],y[46]);
and and3759(ip_58_47,x[58],y[47]);
and and3760(ip_58_48,x[58],y[48]);
and and3761(ip_58_49,x[58],y[49]);
and and3762(ip_58_50,x[58],y[50]);
and and3763(ip_58_51,x[58],y[51]);
and and3764(ip_58_52,x[58],y[52]);
and and3765(ip_58_53,x[58],y[53]);
and and3766(ip_58_54,x[58],y[54]);
and and3767(ip_58_55,x[58],y[55]);
and and3768(ip_58_56,x[58],y[56]);
and and3769(ip_58_57,x[58],y[57]);
and and3770(ip_58_58,x[58],y[58]);
and and3771(ip_58_59,x[58],y[59]);
and and3772(ip_58_60,x[58],y[60]);
and and3773(ip_58_61,x[58],y[61]);
and and3774(ip_58_62,x[58],y[62]);
and and3775(ip_58_63,x[58],y[63]);
and and3776(ip_59_0,x[59],y[0]);
and and3777(ip_59_1,x[59],y[1]);
and and3778(ip_59_2,x[59],y[2]);
and and3779(ip_59_3,x[59],y[3]);
and and3780(ip_59_4,x[59],y[4]);
and and3781(ip_59_5,x[59],y[5]);
and and3782(ip_59_6,x[59],y[6]);
and and3783(ip_59_7,x[59],y[7]);
and and3784(ip_59_8,x[59],y[8]);
and and3785(ip_59_9,x[59],y[9]);
and and3786(ip_59_10,x[59],y[10]);
and and3787(ip_59_11,x[59],y[11]);
and and3788(ip_59_12,x[59],y[12]);
and and3789(ip_59_13,x[59],y[13]);
and and3790(ip_59_14,x[59],y[14]);
and and3791(ip_59_15,x[59],y[15]);
and and3792(ip_59_16,x[59],y[16]);
and and3793(ip_59_17,x[59],y[17]);
and and3794(ip_59_18,x[59],y[18]);
and and3795(ip_59_19,x[59],y[19]);
and and3796(ip_59_20,x[59],y[20]);
and and3797(ip_59_21,x[59],y[21]);
and and3798(ip_59_22,x[59],y[22]);
and and3799(ip_59_23,x[59],y[23]);
and and3800(ip_59_24,x[59],y[24]);
and and3801(ip_59_25,x[59],y[25]);
and and3802(ip_59_26,x[59],y[26]);
and and3803(ip_59_27,x[59],y[27]);
and and3804(ip_59_28,x[59],y[28]);
and and3805(ip_59_29,x[59],y[29]);
and and3806(ip_59_30,x[59],y[30]);
and and3807(ip_59_31,x[59],y[31]);
and and3808(ip_59_32,x[59],y[32]);
and and3809(ip_59_33,x[59],y[33]);
and and3810(ip_59_34,x[59],y[34]);
and and3811(ip_59_35,x[59],y[35]);
and and3812(ip_59_36,x[59],y[36]);
and and3813(ip_59_37,x[59],y[37]);
and and3814(ip_59_38,x[59],y[38]);
and and3815(ip_59_39,x[59],y[39]);
and and3816(ip_59_40,x[59],y[40]);
and and3817(ip_59_41,x[59],y[41]);
and and3818(ip_59_42,x[59],y[42]);
and and3819(ip_59_43,x[59],y[43]);
and and3820(ip_59_44,x[59],y[44]);
and and3821(ip_59_45,x[59],y[45]);
and and3822(ip_59_46,x[59],y[46]);
and and3823(ip_59_47,x[59],y[47]);
and and3824(ip_59_48,x[59],y[48]);
and and3825(ip_59_49,x[59],y[49]);
and and3826(ip_59_50,x[59],y[50]);
and and3827(ip_59_51,x[59],y[51]);
and and3828(ip_59_52,x[59],y[52]);
and and3829(ip_59_53,x[59],y[53]);
and and3830(ip_59_54,x[59],y[54]);
and and3831(ip_59_55,x[59],y[55]);
and and3832(ip_59_56,x[59],y[56]);
and and3833(ip_59_57,x[59],y[57]);
and and3834(ip_59_58,x[59],y[58]);
and and3835(ip_59_59,x[59],y[59]);
and and3836(ip_59_60,x[59],y[60]);
and and3837(ip_59_61,x[59],y[61]);
and and3838(ip_59_62,x[59],y[62]);
and and3839(ip_59_63,x[59],y[63]);
and and3840(ip_60_0,x[60],y[0]);
and and3841(ip_60_1,x[60],y[1]);
and and3842(ip_60_2,x[60],y[2]);
and and3843(ip_60_3,x[60],y[3]);
and and3844(ip_60_4,x[60],y[4]);
and and3845(ip_60_5,x[60],y[5]);
and and3846(ip_60_6,x[60],y[6]);
and and3847(ip_60_7,x[60],y[7]);
and and3848(ip_60_8,x[60],y[8]);
and and3849(ip_60_9,x[60],y[9]);
and and3850(ip_60_10,x[60],y[10]);
and and3851(ip_60_11,x[60],y[11]);
and and3852(ip_60_12,x[60],y[12]);
and and3853(ip_60_13,x[60],y[13]);
and and3854(ip_60_14,x[60],y[14]);
and and3855(ip_60_15,x[60],y[15]);
and and3856(ip_60_16,x[60],y[16]);
and and3857(ip_60_17,x[60],y[17]);
and and3858(ip_60_18,x[60],y[18]);
and and3859(ip_60_19,x[60],y[19]);
and and3860(ip_60_20,x[60],y[20]);
and and3861(ip_60_21,x[60],y[21]);
and and3862(ip_60_22,x[60],y[22]);
and and3863(ip_60_23,x[60],y[23]);
and and3864(ip_60_24,x[60],y[24]);
and and3865(ip_60_25,x[60],y[25]);
and and3866(ip_60_26,x[60],y[26]);
and and3867(ip_60_27,x[60],y[27]);
and and3868(ip_60_28,x[60],y[28]);
and and3869(ip_60_29,x[60],y[29]);
and and3870(ip_60_30,x[60],y[30]);
and and3871(ip_60_31,x[60],y[31]);
and and3872(ip_60_32,x[60],y[32]);
and and3873(ip_60_33,x[60],y[33]);
and and3874(ip_60_34,x[60],y[34]);
and and3875(ip_60_35,x[60],y[35]);
and and3876(ip_60_36,x[60],y[36]);
and and3877(ip_60_37,x[60],y[37]);
and and3878(ip_60_38,x[60],y[38]);
and and3879(ip_60_39,x[60],y[39]);
and and3880(ip_60_40,x[60],y[40]);
and and3881(ip_60_41,x[60],y[41]);
and and3882(ip_60_42,x[60],y[42]);
and and3883(ip_60_43,x[60],y[43]);
and and3884(ip_60_44,x[60],y[44]);
and and3885(ip_60_45,x[60],y[45]);
and and3886(ip_60_46,x[60],y[46]);
and and3887(ip_60_47,x[60],y[47]);
and and3888(ip_60_48,x[60],y[48]);
and and3889(ip_60_49,x[60],y[49]);
and and3890(ip_60_50,x[60],y[50]);
and and3891(ip_60_51,x[60],y[51]);
and and3892(ip_60_52,x[60],y[52]);
and and3893(ip_60_53,x[60],y[53]);
and and3894(ip_60_54,x[60],y[54]);
and and3895(ip_60_55,x[60],y[55]);
and and3896(ip_60_56,x[60],y[56]);
and and3897(ip_60_57,x[60],y[57]);
and and3898(ip_60_58,x[60],y[58]);
and and3899(ip_60_59,x[60],y[59]);
and and3900(ip_60_60,x[60],y[60]);
and and3901(ip_60_61,x[60],y[61]);
and and3902(ip_60_62,x[60],y[62]);
and and3903(ip_60_63,x[60],y[63]);
and and3904(ip_61_0,x[61],y[0]);
and and3905(ip_61_1,x[61],y[1]);
and and3906(ip_61_2,x[61],y[2]);
and and3907(ip_61_3,x[61],y[3]);
and and3908(ip_61_4,x[61],y[4]);
and and3909(ip_61_5,x[61],y[5]);
and and3910(ip_61_6,x[61],y[6]);
and and3911(ip_61_7,x[61],y[7]);
and and3912(ip_61_8,x[61],y[8]);
and and3913(ip_61_9,x[61],y[9]);
and and3914(ip_61_10,x[61],y[10]);
and and3915(ip_61_11,x[61],y[11]);
and and3916(ip_61_12,x[61],y[12]);
and and3917(ip_61_13,x[61],y[13]);
and and3918(ip_61_14,x[61],y[14]);
and and3919(ip_61_15,x[61],y[15]);
and and3920(ip_61_16,x[61],y[16]);
and and3921(ip_61_17,x[61],y[17]);
and and3922(ip_61_18,x[61],y[18]);
and and3923(ip_61_19,x[61],y[19]);
and and3924(ip_61_20,x[61],y[20]);
and and3925(ip_61_21,x[61],y[21]);
and and3926(ip_61_22,x[61],y[22]);
and and3927(ip_61_23,x[61],y[23]);
and and3928(ip_61_24,x[61],y[24]);
and and3929(ip_61_25,x[61],y[25]);
and and3930(ip_61_26,x[61],y[26]);
and and3931(ip_61_27,x[61],y[27]);
and and3932(ip_61_28,x[61],y[28]);
and and3933(ip_61_29,x[61],y[29]);
and and3934(ip_61_30,x[61],y[30]);
and and3935(ip_61_31,x[61],y[31]);
and and3936(ip_61_32,x[61],y[32]);
and and3937(ip_61_33,x[61],y[33]);
and and3938(ip_61_34,x[61],y[34]);
and and3939(ip_61_35,x[61],y[35]);
and and3940(ip_61_36,x[61],y[36]);
and and3941(ip_61_37,x[61],y[37]);
and and3942(ip_61_38,x[61],y[38]);
and and3943(ip_61_39,x[61],y[39]);
and and3944(ip_61_40,x[61],y[40]);
and and3945(ip_61_41,x[61],y[41]);
and and3946(ip_61_42,x[61],y[42]);
and and3947(ip_61_43,x[61],y[43]);
and and3948(ip_61_44,x[61],y[44]);
and and3949(ip_61_45,x[61],y[45]);
and and3950(ip_61_46,x[61],y[46]);
and and3951(ip_61_47,x[61],y[47]);
and and3952(ip_61_48,x[61],y[48]);
and and3953(ip_61_49,x[61],y[49]);
and and3954(ip_61_50,x[61],y[50]);
and and3955(ip_61_51,x[61],y[51]);
and and3956(ip_61_52,x[61],y[52]);
and and3957(ip_61_53,x[61],y[53]);
and and3958(ip_61_54,x[61],y[54]);
and and3959(ip_61_55,x[61],y[55]);
and and3960(ip_61_56,x[61],y[56]);
and and3961(ip_61_57,x[61],y[57]);
and and3962(ip_61_58,x[61],y[58]);
and and3963(ip_61_59,x[61],y[59]);
and and3964(ip_61_60,x[61],y[60]);
and and3965(ip_61_61,x[61],y[61]);
and and3966(ip_61_62,x[61],y[62]);
and and3967(ip_61_63,x[61],y[63]);
and and3968(ip_62_0,x[62],y[0]);
and and3969(ip_62_1,x[62],y[1]);
and and3970(ip_62_2,x[62],y[2]);
and and3971(ip_62_3,x[62],y[3]);
and and3972(ip_62_4,x[62],y[4]);
and and3973(ip_62_5,x[62],y[5]);
and and3974(ip_62_6,x[62],y[6]);
and and3975(ip_62_7,x[62],y[7]);
and and3976(ip_62_8,x[62],y[8]);
and and3977(ip_62_9,x[62],y[9]);
and and3978(ip_62_10,x[62],y[10]);
and and3979(ip_62_11,x[62],y[11]);
and and3980(ip_62_12,x[62],y[12]);
and and3981(ip_62_13,x[62],y[13]);
and and3982(ip_62_14,x[62],y[14]);
and and3983(ip_62_15,x[62],y[15]);
and and3984(ip_62_16,x[62],y[16]);
and and3985(ip_62_17,x[62],y[17]);
and and3986(ip_62_18,x[62],y[18]);
and and3987(ip_62_19,x[62],y[19]);
and and3988(ip_62_20,x[62],y[20]);
and and3989(ip_62_21,x[62],y[21]);
and and3990(ip_62_22,x[62],y[22]);
and and3991(ip_62_23,x[62],y[23]);
and and3992(ip_62_24,x[62],y[24]);
and and3993(ip_62_25,x[62],y[25]);
and and3994(ip_62_26,x[62],y[26]);
and and3995(ip_62_27,x[62],y[27]);
and and3996(ip_62_28,x[62],y[28]);
and and3997(ip_62_29,x[62],y[29]);
and and3998(ip_62_30,x[62],y[30]);
and and3999(ip_62_31,x[62],y[31]);
and and4000(ip_62_32,x[62],y[32]);
and and4001(ip_62_33,x[62],y[33]);
and and4002(ip_62_34,x[62],y[34]);
and and4003(ip_62_35,x[62],y[35]);
and and4004(ip_62_36,x[62],y[36]);
and and4005(ip_62_37,x[62],y[37]);
and and4006(ip_62_38,x[62],y[38]);
and and4007(ip_62_39,x[62],y[39]);
and and4008(ip_62_40,x[62],y[40]);
and and4009(ip_62_41,x[62],y[41]);
and and4010(ip_62_42,x[62],y[42]);
and and4011(ip_62_43,x[62],y[43]);
and and4012(ip_62_44,x[62],y[44]);
and and4013(ip_62_45,x[62],y[45]);
and and4014(ip_62_46,x[62],y[46]);
and and4015(ip_62_47,x[62],y[47]);
and and4016(ip_62_48,x[62],y[48]);
and and4017(ip_62_49,x[62],y[49]);
and and4018(ip_62_50,x[62],y[50]);
and and4019(ip_62_51,x[62],y[51]);
and and4020(ip_62_52,x[62],y[52]);
and and4021(ip_62_53,x[62],y[53]);
and and4022(ip_62_54,x[62],y[54]);
and and4023(ip_62_55,x[62],y[55]);
and and4024(ip_62_56,x[62],y[56]);
and and4025(ip_62_57,x[62],y[57]);
and and4026(ip_62_58,x[62],y[58]);
and and4027(ip_62_59,x[62],y[59]);
and and4028(ip_62_60,x[62],y[60]);
and and4029(ip_62_61,x[62],y[61]);
and and4030(ip_62_62,x[62],y[62]);
and and4031(ip_62_63,x[62],y[63]);
and and4032(ip_63_0,x[63],y[0]);
and and4033(ip_63_1,x[63],y[1]);
and and4034(ip_63_2,x[63],y[2]);
and and4035(ip_63_3,x[63],y[3]);
and and4036(ip_63_4,x[63],y[4]);
and and4037(ip_63_5,x[63],y[5]);
and and4038(ip_63_6,x[63],y[6]);
and and4039(ip_63_7,x[63],y[7]);
and and4040(ip_63_8,x[63],y[8]);
and and4041(ip_63_9,x[63],y[9]);
and and4042(ip_63_10,x[63],y[10]);
and and4043(ip_63_11,x[63],y[11]);
and and4044(ip_63_12,x[63],y[12]);
and and4045(ip_63_13,x[63],y[13]);
and and4046(ip_63_14,x[63],y[14]);
and and4047(ip_63_15,x[63],y[15]);
and and4048(ip_63_16,x[63],y[16]);
and and4049(ip_63_17,x[63],y[17]);
and and4050(ip_63_18,x[63],y[18]);
and and4051(ip_63_19,x[63],y[19]);
and and4052(ip_63_20,x[63],y[20]);
and and4053(ip_63_21,x[63],y[21]);
and and4054(ip_63_22,x[63],y[22]);
and and4055(ip_63_23,x[63],y[23]);
and and4056(ip_63_24,x[63],y[24]);
and and4057(ip_63_25,x[63],y[25]);
and and4058(ip_63_26,x[63],y[26]);
and and4059(ip_63_27,x[63],y[27]);
and and4060(ip_63_28,x[63],y[28]);
and and4061(ip_63_29,x[63],y[29]);
and and4062(ip_63_30,x[63],y[30]);
and and4063(ip_63_31,x[63],y[31]);
and and4064(ip_63_32,x[63],y[32]);
and and4065(ip_63_33,x[63],y[33]);
and and4066(ip_63_34,x[63],y[34]);
and and4067(ip_63_35,x[63],y[35]);
and and4068(ip_63_36,x[63],y[36]);
and and4069(ip_63_37,x[63],y[37]);
and and4070(ip_63_38,x[63],y[38]);
and and4071(ip_63_39,x[63],y[39]);
and and4072(ip_63_40,x[63],y[40]);
and and4073(ip_63_41,x[63],y[41]);
and and4074(ip_63_42,x[63],y[42]);
and and4075(ip_63_43,x[63],y[43]);
and and4076(ip_63_44,x[63],y[44]);
and and4077(ip_63_45,x[63],y[45]);
and and4078(ip_63_46,x[63],y[46]);
and and4079(ip_63_47,x[63],y[47]);
and and4080(ip_63_48,x[63],y[48]);
and and4081(ip_63_49,x[63],y[49]);
and and4082(ip_63_50,x[63],y[50]);
and and4083(ip_63_51,x[63],y[51]);
and and4084(ip_63_52,x[63],y[52]);
and and4085(ip_63_53,x[63],y[53]);
and and4086(ip_63_54,x[63],y[54]);
and and4087(ip_63_55,x[63],y[55]);
and and4088(ip_63_56,x[63],y[56]);
and and4089(ip_63_57,x[63],y[57]);
and and4090(ip_63_58,x[63],y[58]);
and and4091(ip_63_59,x[63],y[59]);
and and4092(ip_63_60,x[63],y[60]);
and and4093(ip_63_61,x[63],y[61]);
and and4094(ip_63_62,x[63],y[62]);
and and4095(ip_63_63,x[63],y[63]);
HA ha0(ip_0_2,ip_1_1,p0,p1);
FA fa0(ip_0_3,ip_1_2,ip_2_1,p2,p3);
FA fa1(ip_3_0,p0,p3,p4,p5);
FA fa2(ip_0_4,ip_1_3,ip_2_2,p6,p7);
FA fa3(ip_3_1,ip_4_0,p7,p8,p9);
FA fa4(p2,p9,p4,p10,p11);
FA fa5(ip_0_5,ip_1_4,ip_2_3,p12,p13);
FA fa6(ip_3_2,ip_4_1,ip_5_0,p14,p15);
FA fa7(p13,p15,p6,p16,p17);
FA fa8(p17,p8,p10,p18,p19);
FA fa9(ip_0_6,ip_1_5,ip_2_4,p20,p21);
FA fa10(ip_3_3,ip_4_2,ip_5_1,p22,p23);
HA ha1(ip_6_0,p21,p24,p25);
FA fa11(p23,p12,p14,p26,p27);
HA ha2(p25,p16,p28,p29);
FA fa12(p27,p29,p18,p30,p31);
FA fa13(ip_0_7,ip_1_6,ip_2_5,p32,p33);
FA fa14(ip_3_4,ip_4_3,ip_5_2,p34,p35);
FA fa15(ip_6_1,ip_7_0,p33,p36,p37);
FA fa16(p35,p20,p22,p38,p39);
FA fa17(p24,p37,p39,p40,p41);
FA fa18(p26,p28,p41,p42,p43);
FA fa19(ip_0_8,ip_1_7,ip_2_6,p44,p45);
FA fa20(ip_3_5,ip_4_4,ip_5_3,p46,p47);
HA ha3(ip_6_2,ip_7_1,p48,p49);
FA fa21(ip_8_0,p49,p45,p50,p51);
HA ha4(p47,p32,p52,p53);
FA fa22(p34,p51,p36,p54,p55);
FA fa23(p53,p55,p38,p56,p57);
FA fa24(p40,p57,p42,p58,p59);
FA fa25(ip_0_9,ip_1_8,ip_2_7,p60,p61);
FA fa26(ip_3_6,ip_4_5,ip_5_4,p62,p63);
HA ha5(ip_6_3,ip_7_2,p64,p65);
FA fa27(ip_8_1,ip_9_0,p48,p66,p67);
FA fa28(p65,p61,p63,p68,p69);
FA fa29(p67,p44,p46,p70,p71);
FA fa30(p50,p52,p69,p72,p73);
FA fa31(p71,p54,p73,p74,p75);
FA fa32(p56,p75,p58,p76,p77);
HA ha6(ip_0_10,ip_1_9,p78,p79);
FA fa33(ip_2_8,ip_3_7,ip_4_6,p80,p81);
HA ha7(ip_5_5,ip_6_4,p82,p83);
HA ha8(ip_7_3,ip_8_2,p84,p85);
FA fa34(ip_9_1,ip_10_0,p64,p86,p87);
FA fa35(p79,p83,p85,p88,p89);
HA ha9(p81,p87,p90,p91);
FA fa36(p60,p62,p66,p92,p93);
HA ha10(p89,p91,p94,p95);
HA ha11(p95,p68,p96,p97);
HA ha12(p93,p70,p98,p99);
FA fa37(p97,p72,p99,p100,p101);
HA ha13(p101,p74,p102,p103);
FA fa38(ip_0_11,ip_1_10,ip_2_9,p104,p105);
HA ha14(ip_3_8,ip_4_7,p106,p107);
FA fa39(ip_5_6,ip_6_5,ip_7_4,p108,p109);
FA fa40(ip_8_3,ip_9_2,ip_10_1,p110,p111);
FA fa41(ip_11_0,p107,p78,p112,p113);
FA fa42(p82,p84,p105,p114,p115);
FA fa43(p109,p111,p113,p116,p117);
FA fa44(p115,p80,p86,p118,p119);
HA ha15(p90,p117,p120,p121);
FA fa45(p88,p94,p119,p122,p123);
HA ha16(p121,p123,p124,p125);
HA ha17(p92,p96,p126,p127);
HA ha18(p125,p127,p128,p129);
FA fa46(p98,p129,p100,p130,p131);
FA fa47(ip_0_12,ip_1_11,ip_2_10,p132,p133);
FA fa48(ip_3_9,ip_4_8,ip_5_7,p134,p135);
HA ha19(ip_6_6,ip_7_5,p136,p137);
FA fa49(ip_8_4,ip_9_3,ip_10_2,p138,p139);
HA ha20(ip_11_1,ip_12_0,p140,p141);
HA ha21(p106,p137,p142,p143);
FA fa50(p141,p133,p135,p144,p145);
FA fa51(p139,p143,p104,p146,p147);
HA ha22(p108,p110,p148,p149);
FA fa52(p112,p114,p145,p150,p151);
FA fa53(p147,p149,p116,p152,p153);
FA fa54(p120,p118,p151,p154,p155);
FA fa55(p153,p122,p124,p156,p157);
HA ha23(p126,p128,p158,p159);
HA ha24(p155,p157,p160,p161);
HA ha25(p159,p161,p162,p163);
HA ha26(ip_0_13,ip_1_12,p164,p165);
FA fa56(ip_2_11,ip_3_10,ip_4_9,p166,p167);
HA ha27(ip_5_8,ip_6_7,p168,p169);
HA ha28(ip_7_6,ip_8_5,p170,p171);
FA fa57(ip_9_4,ip_10_3,ip_11_2,p172,p173);
FA fa58(ip_12_1,ip_13_0,p136,p174,p175);
FA fa59(p140,p165,p169,p176,p177);
FA fa60(p171,p142,p167,p178,p179);
FA fa61(p173,p175,p132,p180,p181);
FA fa62(p134,p138,p177,p182,p183);
FA fa63(p148,p179,p181,p184,p185);
FA fa64(p144,p146,p183,p186,p187);
FA fa65(p185,p150,p152,p188,p189);
FA fa66(p187,p154,p158,p190,p191);
HA ha29(p189,p156,p192,p193);
FA fa67(p160,p162,p191,p194,p195);
HA ha30(ip_0_14,ip_1_13,p196,p197);
HA ha31(ip_2_12,ip_3_11,p198,p199);
FA fa68(ip_4_10,ip_5_9,ip_6_8,p200,p201);
HA ha32(ip_7_7,ip_8_6,p202,p203);
FA fa69(ip_9_5,ip_10_4,ip_11_3,p204,p205);
FA fa70(ip_12_2,ip_13_1,ip_14_0,p206,p207);
HA ha33(p164,p168,p208,p209);
FA fa71(p170,p197,p199,p210,p211);
FA fa72(p203,p201,p205,p212,p213);
FA fa73(p207,p209,p166,p214,p215);
HA ha34(p172,p174,p216,p217);
FA fa74(p211,p176,p213,p218,p219);
HA ha35(p215,p217,p220,p221);
HA ha36(p178,p180,p222,p223);
HA ha37(p221,p182,p224,p225);
HA ha38(p219,p223,p226,p227);
FA fa75(p184,p225,p227,p228,p229);
FA fa76(p186,p229,p188,p230,p231);
FA fa77(p192,p231,p190,p232,p233);
FA fa78(ip_0_15,ip_1_14,ip_2_13,p234,p235);
HA ha39(ip_3_12,ip_4_11,p236,p237);
FA fa79(ip_5_10,ip_6_9,ip_7_8,p238,p239);
FA fa80(ip_8_7,ip_9_6,ip_10_5,p240,p241);
FA fa81(ip_11_4,ip_12_3,ip_13_2,p242,p243);
HA ha40(ip_14_1,ip_15_0,p244,p245);
HA ha41(p196,p198,p246,p247);
HA ha42(p202,p237,p248,p249);
FA fa82(p245,p208,p235,p250,p251);
HA ha43(p239,p241,p252,p253);
FA fa83(p243,p247,p249,p254,p255);
FA fa84(p200,p204,p206,p256,p257);
FA fa85(p253,p210,p216,p258,p259);
FA fa86(p251,p255,p212,p260,p261);
HA ha44(p214,p220,p262,p263);
HA ha45(p257,p222,p264,p265);
FA fa87(p259,p261,p263,p266,p267);
FA fa88(p218,p224,p226,p268,p269);
FA fa89(p265,p267,p269,p270,p271);
HA ha46(p228,p271,p272,p273);
HA ha47(p273,p230,p274,p275);
HA ha48(ip_0_16,ip_1_15,p276,p277);
FA fa90(ip_2_14,ip_3_13,ip_4_12,p278,p279);
FA fa91(ip_5_11,ip_6_10,ip_7_9,p280,p281);
FA fa92(ip_8_8,ip_9_7,ip_10_6,p282,p283);
FA fa93(ip_11_5,ip_12_4,ip_13_3,p284,p285);
FA fa94(ip_14_2,ip_15_1,ip_16_0,p286,p287);
FA fa95(p236,p244,p277,p288,p289);
FA fa96(p246,p248,p279,p290,p291);
HA ha49(p281,p283,p292,p293);
FA fa97(p285,p287,p234,p294,p295);
FA fa98(p238,p240,p242,p296,p297);
HA ha50(p252,p289,p298,p299);
FA fa99(p293,p291,p295,p300,p301);
FA fa100(p299,p250,p254,p302,p303);
FA fa101(p297,p256,p262,p304,p305);
FA fa102(p301,p258,p260,p306,p307);
FA fa103(p264,p303,p305,p308,p309);
FA fa104(p266,p307,p309,p310,p311);
FA fa105(p268,p270,p272,p312,p313);
FA fa106(p311,p274,p313,p314,p315);
HA ha51(ip_0_17,ip_1_16,p316,p317);
FA fa107(ip_2_15,ip_3_14,ip_4_13,p318,p319);
FA fa108(ip_5_12,ip_6_11,ip_7_10,p320,p321);
FA fa109(ip_8_9,ip_9_8,ip_10_7,p322,p323);
FA fa110(ip_11_6,ip_12_5,ip_13_4,p324,p325);
FA fa111(ip_14_3,ip_15_2,ip_16_1,p326,p327);
FA fa112(ip_17_0,p276,p317,p328,p329);
FA fa113(p319,p321,p323,p330,p331);
HA ha52(p325,p327,p332,p333);
FA fa114(p278,p280,p282,p334,p335);
FA fa115(p284,p286,p292,p336,p337);
FA fa116(p329,p333,p288,p338,p339);
HA ha53(p298,p331,p340,p341);
HA ha54(p290,p294,p342,p343);
FA fa117(p335,p337,p339,p344,p345);
FA fa118(p341,p296,p343,p346,p347);
HA ha55(p300,p345,p348,p349);
HA ha56(p302,p347,p350,p351);
HA ha57(p349,p304,p352,p353);
HA ha58(p351,p306,p354,p355);
FA fa119(p308,p353,p355,p356,p357);
FA fa120(p310,p357,p312,p358,p359);
FA fa121(ip_0_18,ip_1_17,ip_2_16,p360,p361);
HA ha59(ip_3_15,ip_4_14,p362,p363);
HA ha60(ip_5_13,ip_6_12,p364,p365);
FA fa122(ip_7_11,ip_8_10,ip_9_9,p366,p367);
HA ha61(ip_10_8,ip_11_7,p368,p369);
FA fa123(ip_12_6,ip_13_5,ip_14_4,p370,p371);
HA ha62(ip_15_3,ip_16_2,p372,p373);
FA fa124(ip_17_1,ip_18_0,p316,p374,p375);
FA fa125(p363,p365,p369,p376,p377);
FA fa126(p373,p361,p367,p378,p379);
FA fa127(p371,p375,p318,p380,p381);
HA ha63(p320,p322,p382,p383);
FA fa128(p324,p326,p332,p384,p385);
FA fa129(p377,p328,p379,p386,p387);
FA fa130(p381,p383,p330,p388,p389);
FA fa131(p340,p385,p334,p390,p391);
FA fa132(p336,p338,p342,p392,p393);
HA ha64(p387,p389,p394,p395);
HA ha65(p391,p395,p396,p397);
FA fa133(p344,p348,p393,p398,p399);
FA fa134(p397,p346,p350,p400,p401);
HA ha66(p352,p399,p402,p403);
FA fa135(p354,p401,p403,p404,p405);
FA fa136(p356,p405,p358,p406,p407);
FA fa137(ip_0_19,ip_1_18,ip_2_17,p408,p409);
HA ha67(ip_3_16,ip_4_15,p410,p411);
FA fa138(ip_5_14,ip_6_13,ip_7_12,p412,p413);
FA fa139(ip_8_11,ip_9_10,ip_10_9,p414,p415);
HA ha68(ip_11_8,ip_12_7,p416,p417);
HA ha69(ip_13_6,ip_14_5,p418,p419);
HA ha70(ip_15_4,ip_16_3,p420,p421);
HA ha71(ip_17_2,ip_18_1,p422,p423);
HA ha72(ip_19_0,p362,p424,p425);
HA ha73(p364,p368,p426,p427);
FA fa140(p372,p411,p417,p428,p429);
FA fa141(p419,p421,p423,p430,p431);
FA fa142(p409,p413,p415,p432,p433);
HA ha74(p425,p427,p434,p435);
HA ha75(p360,p366,p436,p437);
FA fa143(p370,p374,p429,p438,p439);
FA fa144(p431,p435,p376,p440,p441);
HA ha76(p382,p433,p442,p443);
FA fa145(p437,p378,p380,p444,p445);
HA ha77(p439,p441,p446,p447);
FA fa146(p443,p384,p447,p448,p449);
HA ha78(p386,p388,p450,p451);
FA fa147(p394,p445,p390,p452,p453);
HA ha79(p396,p449,p454,p455);
HA ha80(p451,p392,p456,p457);
FA fa148(p453,p455,p457,p458,p459);
FA fa149(p398,p402,p459,p460,p461);
FA fa150(p400,p461,p404,p462,p463);
FA fa151(ip_0_20,ip_1_19,ip_2_18,p464,p465);
FA fa152(ip_3_17,ip_4_16,ip_5_15,p466,p467);
HA ha81(ip_6_14,ip_7_13,p468,p469);
FA fa153(ip_8_12,ip_9_11,ip_10_10,p470,p471);
FA fa154(ip_11_9,ip_12_8,ip_13_7,p472,p473);
FA fa155(ip_14_6,ip_15_5,ip_16_4,p474,p475);
FA fa156(ip_17_3,ip_18_2,ip_19_1,p476,p477);
FA fa157(ip_20_0,p410,p416,p478,p479);
HA ha82(p418,p420,p480,p481);
FA fa158(p422,p469,p424,p482,p483);
HA ha83(p426,p465,p484,p485);
HA ha84(p467,p471,p486,p487);
FA fa159(p473,p475,p477,p488,p489);
FA fa160(p481,p408,p412,p490,p491);
FA fa161(p414,p434,p479,p492,p493);
FA fa162(p483,p485,p487,p494,p495);
FA fa163(p428,p430,p436,p496,p497);
FA fa164(p489,p432,p442,p498,p499);
FA fa165(p491,p493,p495,p500,p501);
HA ha85(p438,p440,p502,p503);
FA fa166(p446,p497,p499,p504,p505);
FA fa167(p501,p503,p444,p506,p507);
FA fa168(p450,p505,p448,p508,p509);
FA fa169(p454,p507,p452,p510,p511);
HA ha86(p456,p509,p512,p513);
FA fa170(p511,p513,p458,p514,p515);
FA fa171(p515,p460,p462,p516,p517);
HA ha87(ip_0_21,ip_1_20,p518,p519);
FA fa172(ip_2_19,ip_3_18,ip_4_17,p520,p521);
FA fa173(ip_5_16,ip_6_15,ip_7_14,p522,p523);
HA ha88(ip_8_13,ip_9_12,p524,p525);
FA fa174(ip_10_11,ip_11_10,ip_12_9,p526,p527);
FA fa175(ip_13_8,ip_14_7,ip_15_6,p528,p529);
FA fa176(ip_16_5,ip_17_4,ip_18_3,p530,p531);
FA fa177(ip_19_2,ip_20_1,ip_21_0,p532,p533);
HA ha89(p468,p519,p534,p535);
FA fa178(p525,p480,p521,p536,p537);
FA fa179(p523,p527,p529,p538,p539);
HA ha90(p531,p533,p540,p541);
FA fa180(p535,p464,p466,p542,p543);
HA ha91(p470,p472,p544,p545);
FA fa181(p474,p476,p484,p546,p547);
FA fa182(p486,p541,p478,p548,p549);
FA fa183(p482,p537,p539,p550,p551);
HA ha92(p545,p488,p552,p553);
FA fa184(p543,p547,p549,p554,p555);
FA fa185(p490,p492,p494,p556,p557);
FA fa186(p551,p553,p496,p558,p559);
HA ha93(p502,p555,p560,p561);
HA ha94(p498,p500,p562,p563);
FA fa187(p557,p559,p561,p564,p565);
HA ha95(p504,p563,p566,p567);
HA ha96(p506,p565,p568,p569);
FA fa188(p567,p508,p512,p570,p571);
FA fa189(p569,p510,p571,p572,p573);
HA ha97(p514,p573,p574,p575);
FA fa190(ip_0_22,ip_1_21,ip_2_20,p576,p577);
HA ha98(ip_3_19,ip_4_18,p578,p579);
HA ha99(ip_5_17,ip_6_16,p580,p581);
FA fa191(ip_7_15,ip_8_14,ip_9_13,p582,p583);
FA fa192(ip_10_12,ip_11_11,ip_12_10,p584,p585);
FA fa193(ip_13_9,ip_14_8,ip_15_7,p586,p587);
FA fa194(ip_16_6,ip_17_5,ip_18_4,p588,p589);
HA ha100(ip_19_3,ip_20_2,p590,p591);
FA fa195(ip_21_1,ip_22_0,p518,p592,p593);
FA fa196(p524,p579,p581,p594,p595);
FA fa197(p591,p534,p577,p596,p597);
HA ha101(p583,p585,p598,p599);
HA ha102(p587,p589,p600,p601);
FA fa198(p593,p520,p522,p602,p603);
HA ha103(p526,p528,p604,p605);
HA ha104(p530,p532,p606,p607);
FA fa199(p540,p595,p599,p608,p609);
FA fa200(p601,p544,p597,p610,p611);
FA fa201(p605,p607,p536,p612,p613);
HA ha105(p538,p603,p614,p615);
FA fa202(p609,p542,p546,p616,p617);
FA fa203(p548,p552,p611,p618,p619);
HA ha106(p613,p615,p620,p621);
FA fa204(p550,p621,p554,p622,p623);
HA ha107(p560,p617,p624,p625);
FA fa205(p619,p556,p558,p626,p627);
FA fa206(p562,p623,p625,p628,p629);
FA fa207(p566,p564,p568,p630,p631);
FA fa208(p627,p629,p631,p632,p633);
HA ha108(p570,p633,p634,p635);
FA fa209(p572,p574,p635,p636,p637);
HA ha109(ip_0_23,ip_1_22,p638,p639);
FA fa210(ip_2_21,ip_3_20,ip_4_19,p640,p641);
FA fa211(ip_5_18,ip_6_17,ip_7_16,p642,p643);
FA fa212(ip_8_15,ip_9_14,ip_10_13,p644,p645);
FA fa213(ip_11_12,ip_12_11,ip_13_10,p646,p647);
FA fa214(ip_14_9,ip_15_8,ip_16_7,p648,p649);
FA fa215(ip_17_6,ip_18_5,ip_19_4,p650,p651);
HA ha110(ip_20_3,ip_21_2,p652,p653);
FA fa216(ip_22_1,ip_23_0,p578,p654,p655);
HA ha111(p580,p590,p656,p657);
FA fa217(p639,p653,p641,p658,p659);
HA ha112(p643,p645,p660,p661);
HA ha113(p647,p649,p662,p663);
FA fa218(p651,p655,p657,p664,p665);
FA fa219(p576,p582,p584,p666,p667);
FA fa220(p586,p588,p592,p668,p669);
FA fa221(p598,p600,p659,p670,p671);
FA fa222(p661,p663,p594,p672,p673);
HA ha114(p604,p606,p674,p675);
FA fa223(p665,p596,p667,p676,p677);
FA fa224(p669,p671,p673,p678,p679);
HA ha115(p675,p602,p680,p681);
FA fa225(p608,p614,p610,p682,p683);
HA ha116(p612,p620,p684,p685);
FA fa226(p677,p679,p681,p686,p687);
FA fa227(p683,p685,p616,p688,p689);
FA fa228(p618,p624,p687,p690,p691);
FA fa229(p622,p689,p691,p692,p693);
FA fa230(p626,p628,p693,p694,p695);
HA ha117(p630,p695,p696,p697);
HA ha118(p632,p634,p698,p699);
FA fa231(p697,p699,p636,p700,p701);
FA fa232(ip_0_24,ip_1_23,ip_2_22,p702,p703);
FA fa233(ip_3_21,ip_4_20,ip_5_19,p704,p705);
FA fa234(ip_6_18,ip_7_17,ip_8_16,p706,p707);
HA ha119(ip_9_15,ip_10_14,p708,p709);
HA ha120(ip_11_13,ip_12_12,p710,p711);
FA fa235(ip_13_11,ip_14_10,ip_15_9,p712,p713);
FA fa236(ip_16_8,ip_17_7,ip_18_6,p714,p715);
HA ha121(ip_19_5,ip_20_4,p716,p717);
HA ha122(ip_21_3,ip_22_2,p718,p719);
HA ha123(ip_23_1,ip_24_0,p720,p721);
FA fa237(p638,p652,p709,p722,p723);
FA fa238(p711,p717,p719,p724,p725);
FA fa239(p721,p656,p703,p726,p727);
HA ha124(p705,p707,p728,p729);
FA fa240(p713,p715,p640,p730,p731);
FA fa241(p642,p644,p646,p732,p733);
FA fa242(p648,p650,p654,p734,p735);
HA ha125(p660,p662,p736,p737);
HA ha126(p723,p725,p738,p739);
FA fa243(p729,p658,p727,p740,p741);
FA fa244(p731,p737,p739,p742,p743);
FA fa245(p664,p674,p733,p744,p745);
HA ha127(p735,p666,p746,p747);
HA ha128(p668,p670,p748,p749);
HA ha129(p672,p741,p750,p751);
HA ha130(p743,p680,p752,p753);
HA ha131(p745,p747,p754,p755);
FA fa246(p749,p751,p676,p756,p757);
FA fa247(p678,p684,p753,p758,p759);
HA ha132(p755,p682,p760,p761);
FA fa248(p757,p686,p759,p762,p763);
FA fa249(p761,p688,p690,p764,p765);
HA ha133(p763,p692,p766,p767);
HA ha134(p765,p767,p768,p769);
FA fa250(p694,p696,p769,p770,p771);
HA ha135(p698,p771,p772,p773);
FA fa251(ip_0_25,ip_1_24,ip_2_23,p774,p775);
FA fa252(ip_3_22,ip_4_21,ip_5_20,p776,p777);
HA ha136(ip_6_19,ip_7_18,p778,p779);
HA ha137(ip_8_17,ip_9_16,p780,p781);
FA fa253(ip_10_15,ip_11_14,ip_12_13,p782,p783);
FA fa254(ip_13_12,ip_14_11,ip_15_10,p784,p785);
FA fa255(ip_16_9,ip_17_8,ip_18_7,p786,p787);
HA ha138(ip_19_6,ip_20_5,p788,p789);
HA ha139(ip_21_4,ip_22_3,p790,p791);
FA fa256(ip_23_2,ip_24_1,ip_25_0,p792,p793);
FA fa257(p708,p710,p716,p794,p795);
FA fa258(p718,p720,p779,p796,p797);
FA fa259(p781,p789,p791,p798,p799);
HA ha140(p775,p777,p800,p801);
FA fa260(p783,p785,p787,p802,p803);
FA fa261(p793,p702,p704,p804,p805);
FA fa262(p706,p712,p714,p806,p807);
FA fa263(p728,p795,p797,p808,p809);
FA fa264(p799,p801,p722,p810,p811);
HA ha141(p724,p736,p812,p813);
FA fa265(p738,p803,p726,p814,p815);
HA ha142(p730,p805,p816,p817);
FA fa266(p807,p809,p811,p818,p819);
FA fa267(p813,p732,p734,p820,p821);
FA fa268(p815,p817,p740,p822,p823);
FA fa269(p742,p746,p748,p824,p825);
HA ha143(p750,p819,p826,p827);
HA ha144(p744,p752,p828,p829);
HA ha145(p754,p821,p830,p831);
FA fa270(p823,p827,p825,p832,p833);
HA ha146(p829,p831,p834,p835);
FA fa271(p756,p760,p833,p836,p837);
FA fa272(p835,p758,p837,p838,p839);
HA ha147(p762,p839,p840,p841);
FA fa273(p764,p766,p841,p842,p843);
FA fa274(p768,p843,p770,p844,p845);
FA fa275(ip_0_26,ip_1_25,ip_2_24,p846,p847);
FA fa276(ip_3_23,ip_4_22,ip_5_21,p848,p849);
FA fa277(ip_6_20,ip_7_19,ip_8_18,p850,p851);
FA fa278(ip_9_17,ip_10_16,ip_11_15,p852,p853);
FA fa279(ip_12_14,ip_13_13,ip_14_12,p854,p855);
FA fa280(ip_15_11,ip_16_10,ip_17_9,p856,p857);
FA fa281(ip_18_8,ip_19_7,ip_20_6,p858,p859);
FA fa282(ip_21_5,ip_22_4,ip_23_3,p860,p861);
FA fa283(ip_24_2,ip_25_1,ip_26_0,p862,p863);
FA fa284(p778,p780,p788,p864,p865);
FA fa285(p790,p847,p849,p866,p867);
HA ha148(p851,p853,p868,p869);
HA ha149(p855,p857,p870,p871);
FA fa286(p859,p861,p863,p872,p873);
FA fa287(p774,p776,p782,p874,p875);
HA ha150(p784,p786,p876,p877);
FA fa288(p792,p800,p865,p878,p879);
HA ha151(p869,p871,p880,p881);
FA fa289(p794,p796,p798,p882,p883);
FA fa290(p867,p873,p877,p884,p885);
FA fa291(p881,p802,p812,p886,p887);
FA fa292(p875,p879,p804,p888,p889);
FA fa293(p806,p808,p810,p890,p891);
HA ha152(p816,p883,p892,p893);
HA ha153(p885,p814,p894,p895);
FA fa294(p887,p889,p893,p896,p897);
FA fa295(p818,p826,p891,p898,p899);
FA fa296(p895,p820,p822,p900,p901);
FA fa297(p828,p830,p897,p902,p903);
FA fa298(p824,p834,p899,p904,p905);
FA fa299(p832,p901,p903,p906,p907);
HA ha154(p905,p836,p908,p909);
FA fa300(p907,p838,p840,p910,p911);
FA fa301(p909,p911,p842,p912,p913);
FA fa302(ip_0_27,ip_1_26,ip_2_25,p914,p915);
FA fa303(ip_3_24,ip_4_23,ip_5_22,p916,p917);
FA fa304(ip_6_21,ip_7_20,ip_8_19,p918,p919);
FA fa305(ip_9_18,ip_10_17,ip_11_16,p920,p921);
HA ha155(ip_12_15,ip_13_14,p922,p923);
HA ha156(ip_14_13,ip_15_12,p924,p925);
HA ha157(ip_16_11,ip_17_10,p926,p927);
HA ha158(ip_18_9,ip_19_8,p928,p929);
FA fa306(ip_20_7,ip_21_6,ip_22_5,p930,p931);
HA ha159(ip_23_4,ip_24_3,p932,p933);
FA fa307(ip_25_2,ip_26_1,ip_27_0,p934,p935);
HA ha160(p923,p925,p936,p937);
FA fa308(p927,p929,p933,p938,p939);
FA fa309(p915,p917,p919,p940,p941);
HA ha161(p921,p931,p942,p943);
HA ha162(p935,p937,p944,p945);
HA ha163(p846,p848,p946,p947);
FA fa310(p850,p852,p854,p948,p949);
FA fa311(p856,p858,p860,p950,p951);
HA ha164(p862,p868,p952,p953);
FA fa312(p870,p939,p943,p954,p955);
HA ha165(p945,p864,p956,p957);
FA fa313(p876,p880,p941,p958,p959);
FA fa314(p947,p953,p866,p960,p961);
FA fa315(p872,p949,p951,p962,p963);
FA fa316(p955,p957,p874,p964,p965);
HA ha166(p878,p959,p966,p967);
FA fa317(p961,p882,p884,p968,p969);
FA fa318(p892,p963,p965,p970,p971);
FA fa319(p967,p886,p888,p972,p973);
HA ha167(p894,p890,p974,p975);
FA fa320(p969,p971,p896,p976,p977);
HA ha168(p973,p975,p978,p979);
HA ha169(p898,p977,p980,p981);
FA fa321(p979,p900,p902,p982,p983);
FA fa322(p981,p904,p906,p984,p985);
HA ha170(p908,p983,p986,p987);
HA ha171(p985,p987,p988,p989);
FA fa323(p989,p910,p912,p990,p991);
FA fa324(ip_0_28,ip_1_27,ip_2_26,p992,p993);
FA fa325(ip_3_25,ip_4_24,ip_5_23,p994,p995);
FA fa326(ip_6_22,ip_7_21,ip_8_20,p996,p997);
HA ha172(ip_9_19,ip_10_18,p998,p999);
HA ha173(ip_11_17,ip_12_16,p1000,p1001);
FA fa327(ip_13_15,ip_14_14,ip_15_13,p1002,p1003);
FA fa328(ip_16_12,ip_17_11,ip_18_10,p1004,p1005);
FA fa329(ip_19_9,ip_20_8,ip_21_7,p1006,p1007);
FA fa330(ip_22_6,ip_23_5,ip_24_4,p1008,p1009);
FA fa331(ip_25_3,ip_26_2,ip_27_1,p1010,p1011);
HA ha174(ip_28_0,p1001,p1012,p1013);
FA fa332(p922,p924,p926,p1014,p1015);
FA fa333(p928,p932,p999,p1016,p1017);
FA fa334(p1003,p1005,p1007,p1018,p1019);
FA fa335(p1009,p1011,p1013,p1020,p1021);
FA fa336(p936,p993,p995,p1022,p1023);
FA fa337(p997,p1015,p1017,p1024,p1025);
HA ha175(p914,p916,p1026,p1027);
FA fa338(p918,p920,p930,p1028,p1029);
FA fa339(p934,p942,p944,p1030,p1031);
FA fa340(p1019,p1021,p1023,p1032,p1033);
FA fa341(p1027,p938,p946,p1034,p1035);
FA fa342(p952,p1025,p1029,p1036,p1037);
HA ha176(p1031,p940,p1038,p1039);
FA fa343(p956,p1033,p1035,p1040,p1041);
FA fa344(p1039,p948,p950,p1042,p1043);
FA fa345(p954,p1037,p958,p1044,p1045);
FA fa346(p960,p966,p1041,p1046,p1047);
FA fa347(p1043,p962,p964,p1048,p1049);
HA ha177(p1045,p1047,p1050,p1051);
HA ha178(p1049,p1051,p1052,p1053);
FA fa348(p968,p970,p974,p1054,p1055);
HA ha179(p1053,p972,p1056,p1057);
FA fa349(p978,p1055,p1057,p1058,p1059);
FA fa350(p976,p980,p1059,p1060,p1061);
FA fa351(p1061,p982,p986,p1062,p1063);
FA fa352(p984,p988,p1063,p1064,p1065);
FA fa353(ip_0_29,ip_1_28,ip_2_27,p1066,p1067);
HA ha180(ip_3_26,ip_4_25,p1068,p1069);
FA fa354(ip_5_24,ip_6_23,ip_7_22,p1070,p1071);
HA ha181(ip_8_21,ip_9_20,p1072,p1073);
HA ha182(ip_10_19,ip_11_18,p1074,p1075);
FA fa355(ip_12_17,ip_13_16,ip_14_15,p1076,p1077);
FA fa356(ip_15_14,ip_16_13,ip_17_12,p1078,p1079);
HA ha183(ip_18_11,ip_19_10,p1080,p1081);
HA ha184(ip_20_9,ip_21_8,p1082,p1083);
HA ha185(ip_22_7,ip_23_6,p1084,p1085);
HA ha186(ip_24_5,ip_25_4,p1086,p1087);
FA fa357(ip_26_3,ip_27_2,ip_28_1,p1088,p1089);
FA fa358(ip_29_0,p1000,p1069,p1090,p1091);
HA ha187(p1073,p1075,p1092,p1093);
FA fa359(p1081,p1083,p1085,p1094,p1095);
FA fa360(p1087,p998,p1012,p1096,p1097);
FA fa361(p1067,p1071,p1077,p1098,p1099);
HA ha188(p1079,p1089,p1100,p1101);
FA fa362(p1093,p1002,p1004,p1102,p1103);
HA ha189(p1006,p1008,p1104,p1105);
FA fa363(p1010,p1091,p1095,p1106,p1107);
FA fa364(p1097,p1101,p992,p1108,p1109);
FA fa365(p994,p996,p1014,p1110,p1111);
HA ha190(p1016,p1026,p1112,p1113);
HA ha191(p1099,p1105,p1114,p1115);
FA fa366(p1018,p1020,p1022,p1116,p1117);
FA fa367(p1103,p1107,p1109,p1118,p1119);
FA fa368(p1111,p1113,p1115,p1120,p1121);
HA ha192(p1024,p1028,p1122,p1123);
FA fa369(p1030,p1038,p1032,p1124,p1125);
HA ha193(p1034,p1117,p1126,p1127);
FA fa370(p1119,p1121,p1123,p1128,p1129);
HA ha194(p1036,p1125,p1130,p1131);
FA fa371(p1127,p1040,p1042,p1132,p1133);
HA ha195(p1129,p1131,p1134,p1135);
HA ha196(p1044,p1046,p1136,p1137);
FA fa372(p1050,p1135,p1048,p1138,p1139);
FA fa373(p1052,p1133,p1137,p1140,p1141);
HA ha197(p1056,p1139,p1142,p1143);
FA fa374(p1054,p1141,p1143,p1144,p1145);
FA fa375(p1058,p1145,p1060,p1146,p1147);
FA fa376(p1147,p1062,p1064,p1148,p1149);
FA fa377(ip_0_30,ip_1_29,ip_2_28,p1150,p1151);
FA fa378(ip_3_27,ip_4_26,ip_5_25,p1152,p1153);
FA fa379(ip_6_24,ip_7_23,ip_8_22,p1154,p1155);
FA fa380(ip_9_21,ip_10_20,ip_11_19,p1156,p1157);
FA fa381(ip_12_18,ip_13_17,ip_14_16,p1158,p1159);
FA fa382(ip_15_15,ip_16_14,ip_17_13,p1160,p1161);
FA fa383(ip_18_12,ip_19_11,ip_20_10,p1162,p1163);
HA ha198(ip_21_9,ip_22_8,p1164,p1165);
FA fa384(ip_23_7,ip_24_6,ip_25_5,p1166,p1167);
FA fa385(ip_26_4,ip_27_3,ip_28_2,p1168,p1169);
FA fa386(ip_29_1,ip_30_0,p1068,p1170,p1171);
HA ha199(p1072,p1074,p1172,p1173);
FA fa387(p1080,p1082,p1084,p1174,p1175);
FA fa388(p1086,p1165,p1092,p1176,p1177);
FA fa389(p1151,p1153,p1155,p1178,p1179);
FA fa390(p1157,p1159,p1161,p1180,p1181);
FA fa391(p1163,p1167,p1169,p1182,p1183);
FA fa392(p1171,p1173,p1066,p1184,p1185);
HA ha200(p1070,p1076,p1186,p1187);
FA fa393(p1078,p1088,p1100,p1188,p1189);
FA fa394(p1175,p1177,p1090,p1190,p1191);
FA fa395(p1094,p1096,p1104,p1192,p1193);
FA fa396(p1179,p1181,p1183,p1194,p1195);
FA fa397(p1185,p1187,p1098,p1196,p1197);
FA fa398(p1112,p1114,p1189,p1198,p1199);
FA fa399(p1191,p1102,p1106,p1200,p1201);
FA fa400(p1108,p1110,p1193,p1202,p1203);
HA ha201(p1195,p1197,p1204,p1205);
HA ha202(p1122,p1199,p1206,p1207);
FA fa401(p1205,p1116,p1118,p1208,p1209);
FA fa402(p1120,p1126,p1201,p1210,p1211);
HA ha203(p1203,p1207,p1212,p1213);
FA fa403(p1124,p1130,p1213,p1214,p1215);
FA fa404(p1128,p1134,p1209,p1216,p1217);
FA fa405(p1211,p1136,p1215,p1218,p1219);
HA ha204(p1132,p1217,p1220,p1221);
HA ha205(p1138,p1142,p1222,p1223);
FA fa406(p1219,p1221,p1140,p1224,p1225);
HA ha206(p1223,p1225,p1226,p1227);
FA fa407(p1144,p1227,p1146,p1228,p1229);
HA ha207(ip_0_31,ip_1_30,p1230,p1231);
HA ha208(ip_2_29,ip_3_28,p1232,p1233);
HA ha209(ip_4_27,ip_5_26,p1234,p1235);
HA ha210(ip_6_25,ip_7_24,p1236,p1237);
FA fa408(ip_8_23,ip_9_22,ip_10_21,p1238,p1239);
FA fa409(ip_11_20,ip_12_19,ip_13_18,p1240,p1241);
FA fa410(ip_14_17,ip_15_16,ip_16_15,p1242,p1243);
FA fa411(ip_17_14,ip_18_13,ip_19_12,p1244,p1245);
HA ha211(ip_20_11,ip_21_10,p1246,p1247);
HA ha212(ip_22_9,ip_23_8,p1248,p1249);
HA ha213(ip_24_7,ip_25_6,p1250,p1251);
FA fa412(ip_26_5,ip_27_4,ip_28_3,p1252,p1253);
FA fa413(ip_29_2,ip_30_1,ip_31_0,p1254,p1255);
HA ha214(p1164,p1231,p1256,p1257);
FA fa414(p1233,p1235,p1237,p1258,p1259);
FA fa415(p1247,p1249,p1251,p1260,p1261);
FA fa416(p1172,p1239,p1241,p1262,p1263);
FA fa417(p1243,p1245,p1253,p1264,p1265);
HA ha215(p1255,p1257,p1266,p1267);
FA fa418(p1150,p1152,p1154,p1268,p1269);
HA ha216(p1156,p1158,p1270,p1271);
HA ha217(p1160,p1162,p1272,p1273);
HA ha218(p1166,p1168,p1274,p1275);
FA fa419(p1170,p1259,p1261,p1276,p1277);
HA ha219(p1267,p1174,p1278,p1279);
FA fa420(p1176,p1186,p1263,p1280,p1281);
FA fa421(p1265,p1271,p1273,p1282,p1283);
HA ha220(p1275,p1178,p1284,p1285);
HA ha221(p1180,p1182,p1286,p1287);
FA fa422(p1184,p1269,p1277,p1288,p1289);
FA fa423(p1279,p1188,p1190,p1290,p1291);
FA fa424(p1281,p1283,p1285,p1292,p1293);
HA ha222(p1287,p1192,p1294,p1295);
FA fa425(p1194,p1196,p1204,p1296,p1297);
HA ha223(p1289,p1198,p1298,p1299);
FA fa426(p1206,p1291,p1293,p1300,p1301);
FA fa427(p1295,p1200,p1202,p1302,p1303);
FA fa428(p1212,p1297,p1299,p1304,p1305);
FA fa429(p1301,p1208,p1210,p1306,p1307);
FA fa430(p1303,p1305,p1214,p1308,p1309);
FA fa431(p1216,p1220,p1307,p1310,p1311);
HA ha224(p1309,p1218,p1312,p1313);
HA ha225(p1222,p1311,p1314,p1315);
HA ha226(p1313,p1224,p1316,p1317);
HA ha227(p1226,p1315,p1318,p1319);
FA fa432(p1317,p1319,p1228,p1320,p1321);
FA fa433(ip_0_32,ip_1_31,ip_2_30,p1322,p1323);
FA fa434(ip_3_29,ip_4_28,ip_5_27,p1324,p1325);
HA ha228(ip_6_26,ip_7_25,p1326,p1327);
FA fa435(ip_8_24,ip_9_23,ip_10_22,p1328,p1329);
HA ha229(ip_11_21,ip_12_20,p1330,p1331);
FA fa436(ip_13_19,ip_14_18,ip_15_17,p1332,p1333);
HA ha230(ip_16_16,ip_17_15,p1334,p1335);
FA fa437(ip_18_14,ip_19_13,ip_20_12,p1336,p1337);
FA fa438(ip_21_11,ip_22_10,ip_23_9,p1338,p1339);
FA fa439(ip_24_8,ip_25_7,ip_26_6,p1340,p1341);
FA fa440(ip_27_5,ip_28_4,ip_29_3,p1342,p1343);
FA fa441(ip_30_2,ip_31_1,ip_32_0,p1344,p1345);
FA fa442(p1230,p1232,p1234,p1346,p1347);
FA fa443(p1236,p1246,p1248,p1348,p1349);
FA fa444(p1250,p1327,p1331,p1350,p1351);
FA fa445(p1335,p1256,p1323,p1352,p1353);
FA fa446(p1325,p1329,p1333,p1354,p1355);
FA fa447(p1337,p1339,p1341,p1356,p1357);
FA fa448(p1343,p1345,p1238,p1358,p1359);
FA fa449(p1240,p1242,p1244,p1360,p1361);
FA fa450(p1252,p1254,p1266,p1362,p1363);
HA ha231(p1347,p1349,p1364,p1365);
FA fa451(p1351,p1258,p1260,p1366,p1367);
HA ha232(p1270,p1272,p1368,p1369);
FA fa452(p1274,p1353,p1355,p1370,p1371);
HA ha233(p1357,p1359,p1372,p1373);
HA ha234(p1365,p1262,p1374,p1375);
HA ha235(p1264,p1278,p1376,p1377);
FA fa453(p1361,p1363,p1369,p1378,p1379);
FA fa454(p1373,p1268,p1276,p1380,p1381);
FA fa455(p1284,p1286,p1367,p1382,p1383);
FA fa456(p1371,p1375,p1377,p1384,p1385);
HA ha236(p1280,p1282,p1386,p1387);
HA ha237(p1379,p1288,p1388,p1389);
FA fa457(p1294,p1381,p1383,p1390,p1391);
FA fa458(p1385,p1387,p1290,p1392,p1393);
FA fa459(p1292,p1298,p1389,p1394,p1395);
FA fa460(p1296,p1391,p1393,p1396,p1397);
FA fa461(p1300,p1395,p1302,p1398,p1399);
HA ha238(p1304,p1397,p1400,p1401);
FA fa462(p1399,p1401,p1306,p1402,p1403);
HA ha239(p1308,p1312,p1404,p1405);
FA fa463(p1403,p1310,p1314,p1406,p1407);
FA fa464(p1405,p1316,p1318,p1408,p1409);
FA fa465(p1407,p1409,p1320,p1410,p1411);
FA fa466(ip_0_33,ip_1_32,ip_2_31,p1412,p1413);
FA fa467(ip_3_30,ip_4_29,ip_5_28,p1414,p1415);
FA fa468(ip_6_27,ip_7_26,ip_8_25,p1416,p1417);
FA fa469(ip_9_24,ip_10_23,ip_11_22,p1418,p1419);
HA ha240(ip_12_21,ip_13_20,p1420,p1421);
FA fa470(ip_14_19,ip_15_18,ip_16_17,p1422,p1423);
HA ha241(ip_17_16,ip_18_15,p1424,p1425);
FA fa471(ip_19_14,ip_20_13,ip_21_12,p1426,p1427);
FA fa472(ip_22_11,ip_23_10,ip_24_9,p1428,p1429);
FA fa473(ip_25_8,ip_26_7,ip_27_6,p1430,p1431);
HA ha242(ip_28_5,ip_29_4,p1432,p1433);
FA fa474(ip_30_3,ip_31_2,ip_32_1,p1434,p1435);
HA ha243(ip_33_0,p1326,p1436,p1437);
FA fa475(p1330,p1334,p1421,p1438,p1439);
FA fa476(p1425,p1433,p1413,p1440,p1441);
FA fa477(p1415,p1417,p1419,p1442,p1443);
HA ha244(p1423,p1427,p1444,p1445);
FA fa478(p1429,p1431,p1435,p1446,p1447);
FA fa479(p1437,p1322,p1324,p1448,p1449);
HA ha245(p1328,p1332,p1450,p1451);
FA fa480(p1336,p1338,p1340,p1452,p1453);
FA fa481(p1342,p1344,p1439,p1454,p1455);
FA fa482(p1441,p1445,p1346,p1456,p1457);
HA ha246(p1348,p1350,p1458,p1459);
HA ha247(p1364,p1443,p1460,p1461);
HA ha248(p1447,p1451,p1462,p1463);
FA fa483(p1352,p1354,p1356,p1464,p1465);
FA fa484(p1358,p1368,p1372,p1466,p1467);
FA fa485(p1449,p1453,p1455,p1468,p1469);
HA ha249(p1457,p1459,p1470,p1471);
FA fa486(p1461,p1463,p1360,p1472,p1473);
FA fa487(p1362,p1374,p1376,p1474,p1475);
HA ha250(p1471,p1366,p1476,p1477);
HA ha251(p1370,p1465,p1478,p1479);
FA fa488(p1467,p1469,p1473,p1480,p1481);
HA ha252(p1378,p1386,p1482,p1483);
FA fa489(p1475,p1477,p1479,p1484,p1485);
FA fa490(p1380,p1382,p1384,p1486,p1487);
FA fa491(p1388,p1481,p1483,p1488,p1489);
FA fa492(p1485,p1390,p1392,p1490,p1491);
FA fa493(p1487,p1489,p1394,p1492,p1493);
HA ha253(p1396,p1400,p1494,p1495);
HA ha254(p1491,p1493,p1496,p1497);
HA ha255(p1398,p1495,p1498,p1499);
FA fa494(p1497,p1499,p1402,p1500,p1501);
FA fa495(p1404,p1501,p1406,p1502,p1503);
HA ha256(p1408,p1503,p1504,p1505);
HA ha257(ip_0_34,ip_1_33,p1506,p1507);
HA ha258(ip_2_32,ip_3_31,p1508,p1509);
FA fa496(ip_4_30,ip_5_29,ip_6_28,p1510,p1511);
FA fa497(ip_7_27,ip_8_26,ip_9_25,p1512,p1513);
FA fa498(ip_10_24,ip_11_23,ip_12_22,p1514,p1515);
HA ha259(ip_13_21,ip_14_20,p1516,p1517);
FA fa499(ip_15_19,ip_16_18,ip_17_17,p1518,p1519);
FA fa500(ip_18_16,ip_19_15,ip_20_14,p1520,p1521);
FA fa501(ip_21_13,ip_22_12,ip_23_11,p1522,p1523);
HA ha260(ip_24_10,ip_25_9,p1524,p1525);
FA fa502(ip_26_8,ip_27_7,ip_28_6,p1526,p1527);
HA ha261(ip_29_5,ip_30_4,p1528,p1529);
HA ha262(ip_31_3,ip_32_2,p1530,p1531);
FA fa503(ip_33_1,ip_34_0,p1420,p1532,p1533);
FA fa504(p1424,p1432,p1507,p1534,p1535);
HA ha263(p1509,p1517,p1536,p1537);
HA ha264(p1525,p1529,p1538,p1539);
FA fa505(p1531,p1436,p1511,p1540,p1541);
FA fa506(p1513,p1515,p1519,p1542,p1543);
HA ha265(p1521,p1523,p1544,p1545);
FA fa507(p1527,p1533,p1537,p1546,p1547);
FA fa508(p1539,p1412,p1414,p1548,p1549);
FA fa509(p1416,p1418,p1422,p1550,p1551);
FA fa510(p1426,p1428,p1430,p1552,p1553);
FA fa511(p1434,p1444,p1535,p1554,p1555);
FA fa512(p1545,p1438,p1440,p1556,p1557);
HA ha266(p1450,p1541,p1558,p1559);
FA fa513(p1543,p1547,p1442,p1560,p1561);
FA fa514(p1446,p1458,p1460,p1562,p1563);
FA fa515(p1462,p1549,p1551,p1564,p1565);
HA ha267(p1553,p1555,p1566,p1567);
HA ha268(p1559,p1448,p1568,p1569);
FA fa516(p1452,p1454,p1456,p1570,p1571);
FA fa517(p1470,p1557,p1561,p1572,p1573);
FA fa518(p1567,p1563,p1565,p1574,p1575);
FA fa519(p1569,p1464,p1466,p1576,p1577);
HA ha269(p1468,p1472,p1578,p1579);
HA ha270(p1476,p1478,p1580,p1581);
FA fa520(p1571,p1573,p1474,p1582,p1583);
HA ha271(p1482,p1575,p1584,p1585);
HA ha272(p1579,p1581,p1586,p1587);
FA fa521(p1480,p1577,p1583,p1588,p1589);
FA fa522(p1585,p1587,p1484,p1590,p1591);
FA fa523(p1486,p1488,p1589,p1592,p1593);
FA fa524(p1591,p1490,p1492,p1594,p1595);
FA fa525(p1494,p1496,p1593,p1596,p1597);
HA ha273(p1498,p1595,p1598,p1599);
HA ha274(p1597,p1599,p1600,p1601);
FA fa526(p1500,p1601,p1502,p1602,p1603);
FA fa527(ip_0_35,ip_1_34,ip_2_33,p1604,p1605);
FA fa528(ip_3_32,ip_4_31,ip_5_30,p1606,p1607);
FA fa529(ip_6_29,ip_7_28,ip_8_27,p1608,p1609);
FA fa530(ip_9_26,ip_10_25,ip_11_24,p1610,p1611);
FA fa531(ip_12_23,ip_13_22,ip_14_21,p1612,p1613);
FA fa532(ip_15_20,ip_16_19,ip_17_18,p1614,p1615);
FA fa533(ip_18_17,ip_19_16,ip_20_15,p1616,p1617);
FA fa534(ip_21_14,ip_22_13,ip_23_12,p1618,p1619);
HA ha275(ip_24_11,ip_25_10,p1620,p1621);
HA ha276(ip_26_9,ip_27_8,p1622,p1623);
FA fa535(ip_28_7,ip_29_6,ip_30_5,p1624,p1625);
FA fa536(ip_31_4,ip_32_3,ip_33_2,p1626,p1627);
FA fa537(ip_34_1,ip_35_0,p1506,p1628,p1629);
FA fa538(p1508,p1516,p1524,p1630,p1631);
HA ha277(p1528,p1530,p1632,p1633);
FA fa539(p1621,p1623,p1536,p1634,p1635);
FA fa540(p1538,p1605,p1607,p1636,p1637);
FA fa541(p1609,p1611,p1613,p1638,p1639);
FA fa542(p1615,p1617,p1619,p1640,p1641);
FA fa543(p1625,p1627,p1629,p1642,p1643);
HA ha278(p1633,p1510,p1644,p1645);
FA fa544(p1512,p1514,p1518,p1646,p1647);
HA ha279(p1520,p1522,p1648,p1649);
HA ha280(p1526,p1532,p1650,p1651);
HA ha281(p1544,p1631,p1652,p1653);
HA ha282(p1635,p1534,p1654,p1655);
FA fa545(p1637,p1639,p1641,p1656,p1657);
FA fa546(p1643,p1645,p1649,p1658,p1659);
FA fa547(p1651,p1653,p1540,p1660,p1661);
HA ha283(p1542,p1546,p1662,p1663);
HA ha284(p1558,p1647,p1664,p1665);
FA fa548(p1655,p1548,p1550,p1666,p1667);
FA fa549(p1552,p1554,p1566,p1668,p1669);
FA fa550(p1657,p1659,p1661,p1670,p1671);
FA fa551(p1663,p1665,p1556,p1672,p1673);
FA fa552(p1560,p1568,p1562,p1674,p1675);
HA ha285(p1564,p1667,p1676,p1677);
FA fa553(p1669,p1671,p1673,p1678,p1679);
FA fa554(p1570,p1572,p1578,p1680,p1681);
HA ha286(p1580,p1675,p1682,p1683);
FA fa555(p1677,p1574,p1584,p1684,p1685);
FA fa556(p1586,p1679,p1683,p1686,p1687);
HA ha287(p1576,p1582,p1688,p1689);
HA ha288(p1681,p1685,p1690,p1691);
HA ha289(p1687,p1689,p1692,p1693);
HA ha290(p1588,p1590,p1694,p1695);
FA fa557(p1691,p1693,p1695,p1696,p1697);
HA ha291(p1592,p1697,p1698,p1699);
HA ha292(p1699,p1594,p1700,p1701);
FA fa558(p1596,p1598,p1600,p1702,p1703);
HA ha293(p1701,p1703,p1704,p1705);
FA fa559(ip_0_36,ip_1_35,ip_2_34,p1706,p1707);
FA fa560(ip_3_33,ip_4_32,ip_5_31,p1708,p1709);
FA fa561(ip_6_30,ip_7_29,ip_8_28,p1710,p1711);
HA ha294(ip_9_27,ip_10_26,p1712,p1713);
HA ha295(ip_11_25,ip_12_24,p1714,p1715);
FA fa562(ip_13_23,ip_14_22,ip_15_21,p1716,p1717);
HA ha296(ip_16_20,ip_17_19,p1718,p1719);
FA fa563(ip_18_18,ip_19_17,ip_20_16,p1720,p1721);
FA fa564(ip_21_15,ip_22_14,ip_23_13,p1722,p1723);
FA fa565(ip_24_12,ip_25_11,ip_26_10,p1724,p1725);
HA ha297(ip_27_9,ip_28_8,p1726,p1727);
HA ha298(ip_29_7,ip_30_6,p1728,p1729);
FA fa566(ip_31_5,ip_32_4,ip_33_3,p1730,p1731);
FA fa567(ip_34_2,ip_35_1,ip_36_0,p1732,p1733);
HA ha299(p1620,p1622,p1734,p1735);
FA fa568(p1713,p1715,p1719,p1736,p1737);
HA ha300(p1727,p1729,p1738,p1739);
FA fa569(p1632,p1707,p1709,p1740,p1741);
HA ha301(p1711,p1717,p1742,p1743);
FA fa570(p1721,p1723,p1725,p1744,p1745);
FA fa571(p1731,p1733,p1735,p1746,p1747);
FA fa572(p1739,p1604,p1606,p1748,p1749);
HA ha302(p1608,p1610,p1750,p1751);
FA fa573(p1612,p1614,p1616,p1752,p1753);
HA ha303(p1618,p1624,p1754,p1755);
HA ha304(p1626,p1628,p1756,p1757);
HA ha305(p1737,p1743,p1758,p1759);
HA ha306(p1630,p1634,p1760,p1761);
FA fa574(p1644,p1648,p1650,p1762,p1763);
FA fa575(p1652,p1741,p1745,p1764,p1765);
FA fa576(p1747,p1751,p1755,p1766,p1767);
FA fa577(p1757,p1759,p1636,p1768,p1769);
HA ha307(p1638,p1640,p1770,p1771);
FA fa578(p1642,p1654,p1749,p1772,p1773);
FA fa579(p1753,p1761,p1646,p1774,p1775);
FA fa580(p1662,p1664,p1763,p1776,p1777);
FA fa581(p1765,p1767,p1769,p1778,p1779);
FA fa582(p1771,p1656,p1658,p1780,p1781);
HA ha308(p1660,p1773,p1782,p1783);
FA fa583(p1775,p1777,p1779,p1784,p1785);
HA ha309(p1783,p1666,p1786,p1787);
HA ha310(p1668,p1670,p1788,p1789);
FA fa584(p1672,p1676,p1781,p1790,p1791);
FA fa585(p1674,p1682,p1785,p1792,p1793);
FA fa586(p1787,p1789,p1678,p1794,p1795);
FA fa587(p1791,p1680,p1688,p1796,p1797);
FA fa588(p1793,p1795,p1684,p1798,p1799);
FA fa589(p1686,p1690,p1692,p1800,p1801);
HA ha311(p1694,p1797,p1802,p1803);
FA fa590(p1799,p1801,p1803,p1804,p1805);
FA fa591(p1696,p1698,p1805,p1806,p1807);
FA fa592(p1700,p1807,p1702,p1808,p1809);
FA fa593(ip_0_37,ip_1_36,ip_2_35,p1810,p1811);
FA fa594(ip_3_34,ip_4_33,ip_5_32,p1812,p1813);
FA fa595(ip_6_31,ip_7_30,ip_8_29,p1814,p1815);
FA fa596(ip_9_28,ip_10_27,ip_11_26,p1816,p1817);
FA fa597(ip_12_25,ip_13_24,ip_14_23,p1818,p1819);
FA fa598(ip_15_22,ip_16_21,ip_17_20,p1820,p1821);
HA ha312(ip_18_19,ip_19_18,p1822,p1823);
HA ha313(ip_20_17,ip_21_16,p1824,p1825);
FA fa599(ip_22_15,ip_23_14,ip_24_13,p1826,p1827);
HA ha314(ip_25_12,ip_26_11,p1828,p1829);
FA fa600(ip_27_10,ip_28_9,ip_29_8,p1830,p1831);
FA fa601(ip_30_7,ip_31_6,ip_32_5,p1832,p1833);
FA fa602(ip_33_4,ip_34_3,ip_35_2,p1834,p1835);
FA fa603(ip_36_1,ip_37_0,p1712,p1836,p1837);
FA fa604(p1714,p1718,p1726,p1838,p1839);
HA ha315(p1728,p1823,p1840,p1841);
HA ha316(p1825,p1829,p1842,p1843);
FA fa605(p1734,p1738,p1811,p1844,p1845);
FA fa606(p1813,p1815,p1817,p1846,p1847);
FA fa607(p1819,p1821,p1827,p1848,p1849);
FA fa608(p1831,p1833,p1835,p1850,p1851);
FA fa609(p1837,p1841,p1843,p1852,p1853);
FA fa610(p1706,p1708,p1710,p1854,p1855);
HA ha317(p1716,p1720,p1856,p1857);
HA ha318(p1722,p1724,p1858,p1859);
FA fa611(p1730,p1732,p1742,p1860,p1861);
FA fa612(p1839,p1736,p1750,p1862,p1863);
FA fa613(p1754,p1756,p1758,p1864,p1865);
FA fa614(p1845,p1847,p1849,p1866,p1867);
HA ha319(p1851,p1853,p1868,p1869);
HA ha320(p1857,p1859,p1870,p1871);
FA fa615(p1740,p1744,p1746,p1872,p1873);
FA fa616(p1760,p1855,p1861,p1874,p1875);
HA ha321(p1869,p1871,p1876,p1877);
HA ha322(p1748,p1752,p1878,p1879);
FA fa617(p1770,p1863,p1865,p1880,p1881);
FA fa618(p1867,p1877,p1762,p1882,p1883);
FA fa619(p1764,p1766,p1768,p1884,p1885);
FA fa620(p1873,p1875,p1879,p1886,p1887);
FA fa621(p1772,p1774,p1782,p1888,p1889);
HA ha323(p1881,p1883,p1890,p1891);
FA fa622(p1776,p1778,p1885,p1892,p1893);
FA fa623(p1887,p1891,p1780,p1894,p1895);
HA ha324(p1786,p1788,p1896,p1897);
FA fa624(p1889,p1784,p1893,p1898,p1899);
FA fa625(p1895,p1897,p1790,p1900,p1901);
FA fa626(p1792,p1794,p1899,p1902,p1903);
FA fa627(p1901,p1796,p1798,p1904,p1905);
FA fa628(p1802,p1903,p1800,p1906,p1907);
HA ha325(p1905,p1907,p1908,p1909);
FA fa629(p1804,p1909,p1806,p1910,p1911);
FA fa630(ip_0_38,ip_1_37,ip_2_36,p1912,p1913);
FA fa631(ip_3_35,ip_4_34,ip_5_33,p1914,p1915);
FA fa632(ip_6_32,ip_7_31,ip_8_30,p1916,p1917);
FA fa633(ip_9_29,ip_10_28,ip_11_27,p1918,p1919);
FA fa634(ip_12_26,ip_13_25,ip_14_24,p1920,p1921);
FA fa635(ip_15_23,ip_16_22,ip_17_21,p1922,p1923);
HA ha326(ip_18_20,ip_19_19,p1924,p1925);
HA ha327(ip_20_18,ip_21_17,p1926,p1927);
FA fa636(ip_22_16,ip_23_15,ip_24_14,p1928,p1929);
FA fa637(ip_25_13,ip_26_12,ip_27_11,p1930,p1931);
HA ha328(ip_28_10,ip_29_9,p1932,p1933);
FA fa638(ip_30_8,ip_31_7,ip_32_6,p1934,p1935);
FA fa639(ip_33_5,ip_34_4,ip_35_3,p1936,p1937);
HA ha329(ip_36_2,ip_37_1,p1938,p1939);
HA ha330(ip_38_0,p1822,p1940,p1941);
FA fa640(p1824,p1828,p1925,p1942,p1943);
FA fa641(p1927,p1933,p1939,p1944,p1945);
FA fa642(p1840,p1842,p1913,p1946,p1947);
FA fa643(p1915,p1917,p1919,p1948,p1949);
FA fa644(p1921,p1923,p1929,p1950,p1951);
HA ha331(p1931,p1935,p1952,p1953);
FA fa645(p1937,p1941,p1810,p1954,p1955);
FA fa646(p1812,p1814,p1816,p1956,p1957);
HA ha332(p1818,p1820,p1958,p1959);
FA fa647(p1826,p1830,p1832,p1960,p1961);
HA ha333(p1834,p1836,p1962,p1963);
FA fa648(p1943,p1945,p1953,p1964,p1965);
HA ha334(p1838,p1856,p1966,p1967);
HA ha335(p1858,p1947,p1968,p1969);
FA fa649(p1949,p1951,p1955,p1970,p1971);
HA ha336(p1959,p1963,p1972,p1973);
FA fa650(p1844,p1846,p1848,p1974,p1975);
FA fa651(p1850,p1852,p1868,p1976,p1977);
FA fa652(p1870,p1957,p1961,p1978,p1979);
FA fa653(p1965,p1967,p1969,p1980,p1981);
HA ha337(p1973,p1854,p1982,p1983);
FA fa654(p1860,p1876,p1971,p1984,p1985);
HA ha338(p1862,p1864,p1986,p1987);
HA ha339(p1866,p1878,p1988,p1989);
FA fa655(p1975,p1977,p1979,p1990,p1991);
HA ha340(p1981,p1983,p1992,p1993);
FA fa656(p1872,p1874,p1985,p1994,p1995);
FA fa657(p1987,p1989,p1993,p1996,p1997);
HA ha341(p1880,p1882,p1998,p1999);
FA fa658(p1890,p1991,p1884,p2000,p2001);
FA fa659(p1886,p1995,p1997,p2002,p2003);
FA fa660(p1999,p1888,p1896,p2004,p2005);
FA fa661(p2001,p1892,p1894,p2006,p2007);
FA fa662(p2003,p2005,p1898,p2008,p2009);
FA fa663(p1900,p2007,p2009,p2010,p2011);
FA fa664(p1902,p2011,p1904,p2012,p2013);
HA ha342(p1906,p1908,p2014,p2015);
FA fa665(p2013,p2015,p1910,p2016,p2017);
FA fa666(ip_0_39,ip_1_38,ip_2_37,p2018,p2019);
HA ha343(ip_3_36,ip_4_35,p2020,p2021);
HA ha344(ip_5_34,ip_6_33,p2022,p2023);
FA fa667(ip_7_32,ip_8_31,ip_9_30,p2024,p2025);
FA fa668(ip_10_29,ip_11_28,ip_12_27,p2026,p2027);
FA fa669(ip_13_26,ip_14_25,ip_15_24,p2028,p2029);
HA ha345(ip_16_23,ip_17_22,p2030,p2031);
FA fa670(ip_18_21,ip_19_20,ip_20_19,p2032,p2033);
HA ha346(ip_21_18,ip_22_17,p2034,p2035);
FA fa671(ip_23_16,ip_24_15,ip_25_14,p2036,p2037);
HA ha347(ip_26_13,ip_27_12,p2038,p2039);
FA fa672(ip_28_11,ip_29_10,ip_30_9,p2040,p2041);
FA fa673(ip_31_8,ip_32_7,ip_33_6,p2042,p2043);
FA fa674(ip_34_5,ip_35_4,ip_36_3,p2044,p2045);
FA fa675(ip_37_2,ip_38_1,ip_39_0,p2046,p2047);
HA ha348(p1924,p1926,p2048,p2049);
FA fa676(p1932,p1938,p2021,p2050,p2051);
HA ha349(p2023,p2031,p2052,p2053);
FA fa677(p2035,p2039,p1940,p2054,p2055);
FA fa678(p2019,p2025,p2027,p2056,p2057);
FA fa679(p2029,p2033,p2037,p2058,p2059);
HA ha350(p2041,p2043,p2060,p2061);
FA fa680(p2045,p2047,p2049,p2062,p2063);
FA fa681(p2053,p1912,p1914,p2064,p2065);
FA fa682(p1916,p1918,p1920,p2066,p2067);
FA fa683(p1922,p1928,p1930,p2068,p2069);
HA ha351(p1934,p1936,p2070,p2071);
HA ha352(p1952,p2051,p2072,p2073);
FA fa684(p2055,p2061,p1942,p2074,p2075);
HA ha353(p1944,p1958,p2076,p2077);
FA fa685(p1962,p2057,p2059,p2078,p2079);
FA fa686(p2063,p2071,p2073,p2080,p2081);
FA fa687(p1946,p1948,p1950,p2082,p2083);
HA ha354(p1954,p1966,p2084,p2085);
HA ha355(p1968,p1972,p2086,p2087);
FA fa688(p2065,p2067,p2069,p2088,p2089);
FA fa689(p2075,p2077,p1956,p2090,p2091);
FA fa690(p1960,p1964,p2079,p2092,p2093);
FA fa691(p2081,p2085,p2087,p2094,p2095);
HA ha356(p1970,p1982,p2096,p2097);
FA fa692(p2083,p2089,p2091,p2098,p2099);
HA ha357(p1974,p1976,p2100,p2101);
FA fa693(p1978,p1980,p1986,p2102,p2103);
FA fa694(p1988,p1992,p2093,p2104,p2105);
FA fa695(p2095,p2097,p1984,p2106,p2107);
FA fa696(p2099,p2101,p1990,p2108,p2109);
FA fa697(p1998,p2103,p2105,p2110,p2111);
FA fa698(p2107,p1994,p1996,p2112,p2113);
FA fa699(p2109,p2000,p2111,p2114,p2115);
HA ha358(p2002,p2113,p2116,p2117);
FA fa700(p2004,p2115,p2117,p2118,p2119);
FA fa701(p2006,p2008,p2119,p2120,p2121);
FA fa702(p2010,p2121,p2014,p2122,p2123);
HA ha359(p2012,p2123,p2124,p2125);
HA ha360(ip_0_40,ip_1_39,p2126,p2127);
HA ha361(ip_2_38,ip_3_37,p2128,p2129);
FA fa703(ip_4_36,ip_5_35,ip_6_34,p2130,p2131);
FA fa704(ip_7_33,ip_8_32,ip_9_31,p2132,p2133);
HA ha362(ip_10_30,ip_11_29,p2134,p2135);
FA fa705(ip_12_28,ip_13_27,ip_14_26,p2136,p2137);
HA ha363(ip_15_25,ip_16_24,p2138,p2139);
FA fa706(ip_17_23,ip_18_22,ip_19_21,p2140,p2141);
FA fa707(ip_20_20,ip_21_19,ip_22_18,p2142,p2143);
FA fa708(ip_23_17,ip_24_16,ip_25_15,p2144,p2145);
HA ha364(ip_26_14,ip_27_13,p2146,p2147);
FA fa709(ip_28_12,ip_29_11,ip_30_10,p2148,p2149);
HA ha365(ip_31_9,ip_32_8,p2150,p2151);
HA ha366(ip_33_7,ip_34_6,p2152,p2153);
FA fa710(ip_35_5,ip_36_4,ip_37_3,p2154,p2155);
HA ha367(ip_38_2,ip_39_1,p2156,p2157);
FA fa711(ip_40_0,p2020,p2022,p2158,p2159);
FA fa712(p2030,p2034,p2038,p2160,p2161);
HA ha368(p2127,p2129,p2162,p2163);
FA fa713(p2135,p2139,p2147,p2164,p2165);
HA ha369(p2151,p2153,p2166,p2167);
FA fa714(p2157,p2048,p2052,p2168,p2169);
FA fa715(p2131,p2133,p2137,p2170,p2171);
FA fa716(p2141,p2143,p2145,p2172,p2173);
FA fa717(p2149,p2155,p2163,p2174,p2175);
FA fa718(p2167,p2018,p2024,p2176,p2177);
HA ha370(p2026,p2028,p2178,p2179);
HA ha371(p2032,p2036,p2180,p2181);
FA fa719(p2040,p2042,p2044,p2182,p2183);
HA ha372(p2046,p2060,p2184,p2185);
FA fa720(p2159,p2161,p2165,p2186,p2187);
FA fa721(p2050,p2054,p2070,p2188,p2189);
HA ha373(p2072,p2169,p2190,p2191);
FA fa722(p2171,p2173,p2175,p2192,p2193);
FA fa723(p2179,p2181,p2185,p2194,p2195);
FA fa724(p2056,p2058,p2062,p2196,p2197);
HA ha374(p2076,p2177,p2198,p2199);
FA fa725(p2183,p2187,p2191,p2200,p2201);
FA fa726(p2064,p2066,p2068,p2202,p2203);
FA fa727(p2074,p2084,p2086,p2204,p2205);
HA ha375(p2189,p2193,p2206,p2207);
HA ha376(p2195,p2199,p2208,p2209);
FA fa728(p2078,p2080,p2197,p2210,p2211);
FA fa729(p2201,p2207,p2209,p2212,p2213);
FA fa730(p2082,p2088,p2090,p2214,p2215);
HA ha377(p2096,p2203,p2216,p2217);
HA ha378(p2205,p2092,p2218,p2219);
FA fa731(p2094,p2100,p2211,p2220,p2221);
FA fa732(p2213,p2217,p2098,p2222,p2223);
FA fa733(p2215,p2219,p2102,p2224,p2225);
HA ha379(p2104,p2106,p2226,p2227);
HA ha380(p2221,p2223,p2228,p2229);
HA ha381(p2108,p2225,p2230,p2231);
FA fa734(p2227,p2229,p2110,p2232,p2233);
FA fa735(p2231,p2112,p2116,p2234,p2235);
FA fa736(p2233,p2114,p2235,p2236,p2237);
FA fa737(p2118,p2237,p2120,p2238,p2239);
FA fa738(p2239,p2122,p2124,p2240,p2241);
FA fa739(ip_0_41,ip_1_40,ip_2_39,p2242,p2243);
FA fa740(ip_3_38,ip_4_37,ip_5_36,p2244,p2245);
HA ha382(ip_6_35,ip_7_34,p2246,p2247);
HA ha383(ip_8_33,ip_9_32,p2248,p2249);
FA fa741(ip_10_31,ip_11_30,ip_12_29,p2250,p2251);
HA ha384(ip_13_28,ip_14_27,p2252,p2253);
FA fa742(ip_15_26,ip_16_25,ip_17_24,p2254,p2255);
HA ha385(ip_18_23,ip_19_22,p2256,p2257);
HA ha386(ip_20_21,ip_21_20,p2258,p2259);
HA ha387(ip_22_19,ip_23_18,p2260,p2261);
FA fa743(ip_24_17,ip_25_16,ip_26_15,p2262,p2263);
HA ha388(ip_27_14,ip_28_13,p2264,p2265);
HA ha389(ip_29_12,ip_30_11,p2266,p2267);
FA fa744(ip_31_10,ip_32_9,ip_33_8,p2268,p2269);
FA fa745(ip_34_7,ip_35_6,ip_36_5,p2270,p2271);
HA ha390(ip_37_4,ip_38_3,p2272,p2273);
FA fa746(ip_39_2,ip_40_1,ip_41_0,p2274,p2275);
FA fa747(p2126,p2128,p2134,p2276,p2277);
HA ha391(p2138,p2146,p2278,p2279);
HA ha392(p2150,p2152,p2280,p2281);
FA fa748(p2156,p2247,p2249,p2282,p2283);
FA fa749(p2253,p2257,p2259,p2284,p2285);
HA ha393(p2261,p2265,p2286,p2287);
HA ha394(p2267,p2273,p2288,p2289);
FA fa750(p2162,p2166,p2243,p2290,p2291);
FA fa751(p2245,p2251,p2255,p2292,p2293);
FA fa752(p2263,p2269,p2271,p2294,p2295);
HA ha395(p2275,p2279,p2296,p2297);
HA ha396(p2281,p2287,p2298,p2299);
HA ha397(p2289,p2130,p2300,p2301);
HA ha398(p2132,p2136,p2302,p2303);
FA fa753(p2140,p2142,p2144,p2304,p2305);
FA fa754(p2148,p2154,p2277,p2306,p2307);
FA fa755(p2283,p2285,p2297,p2308,p2309);
HA ha399(p2299,p2158,p2310,p2311);
FA fa756(p2160,p2164,p2178,p2312,p2313);
FA fa757(p2180,p2184,p2291,p2314,p2315);
HA ha400(p2293,p2295,p2316,p2317);
FA fa758(p2301,p2303,p2168,p2318,p2319);
FA fa759(p2170,p2172,p2174,p2320,p2321);
HA ha401(p2190,p2305,p2322,p2323);
FA fa760(p2307,p2309,p2311,p2324,p2325);
FA fa761(p2317,p2176,p2182,p2326,p2327);
FA fa762(p2186,p2198,p2313,p2328,p2329);
FA fa763(p2315,p2319,p2323,p2330,p2331);
FA fa764(p2188,p2192,p2194,p2332,p2333);
FA fa765(p2206,p2208,p2321,p2334,p2335);
FA fa766(p2325,p2196,p2200,p2336,p2337);
FA fa767(p2327,p2329,p2331,p2338,p2339);
FA fa768(p2202,p2204,p2216,p2340,p2341);
FA fa769(p2333,p2335,p2210,p2342,p2343);
FA fa770(p2212,p2218,p2337,p2344,p2345);
FA fa771(p2339,p2214,p2341,p2346,p2347);
FA fa772(p2343,p2220,p2222,p2348,p2349);
HA ha402(p2226,p2228,p2350,p2351);
HA ha403(p2345,p2224,p2352,p2353);
HA ha404(p2230,p2347,p2354,p2355);
FA fa773(p2351,p2349,p2353,p2356,p2357);
FA fa774(p2355,p2232,p2357,p2358,p2359);
HA ha405(p2234,p2359,p2360,p2361);
FA fa775(p2236,p2361,p2238,p2362,p2363);
HA ha406(ip_0_42,ip_1_41,p2364,p2365);
HA ha407(ip_2_40,ip_3_39,p2366,p2367);
FA fa776(ip_4_38,ip_5_37,ip_6_36,p2368,p2369);
HA ha408(ip_7_35,ip_8_34,p2370,p2371);
FA fa777(ip_9_33,ip_10_32,ip_11_31,p2372,p2373);
FA fa778(ip_12_30,ip_13_29,ip_14_28,p2374,p2375);
FA fa779(ip_15_27,ip_16_26,ip_17_25,p2376,p2377);
FA fa780(ip_18_24,ip_19_23,ip_20_22,p2378,p2379);
FA fa781(ip_21_21,ip_22_20,ip_23_19,p2380,p2381);
HA ha409(ip_24_18,ip_25_17,p2382,p2383);
FA fa782(ip_26_16,ip_27_15,ip_28_14,p2384,p2385);
FA fa783(ip_29_13,ip_30_12,ip_31_11,p2386,p2387);
FA fa784(ip_32_10,ip_33_9,ip_34_8,p2388,p2389);
HA ha410(ip_35_7,ip_36_6,p2390,p2391);
FA fa785(ip_37_5,ip_38_4,ip_39_3,p2392,p2393);
FA fa786(ip_40_2,ip_41_1,ip_42_0,p2394,p2395);
FA fa787(p2246,p2248,p2252,p2396,p2397);
FA fa788(p2256,p2258,p2260,p2398,p2399);
HA ha411(p2264,p2266,p2400,p2401);
FA fa789(p2272,p2365,p2367,p2402,p2403);
FA fa790(p2371,p2383,p2391,p2404,p2405);
HA ha412(p2278,p2280,p2406,p2407);
HA ha413(p2286,p2288,p2408,p2409);
FA fa791(p2369,p2373,p2375,p2410,p2411);
FA fa792(p2377,p2379,p2381,p2412,p2413);
HA ha414(p2385,p2387,p2414,p2415);
HA ha415(p2389,p2393,p2416,p2417);
HA ha416(p2395,p2401,p2418,p2419);
FA fa793(p2242,p2244,p2250,p2420,p2421);
HA ha417(p2254,p2262,p2422,p2423);
HA ha418(p2268,p2270,p2424,p2425);
FA fa794(p2274,p2296,p2298,p2426,p2427);
FA fa795(p2397,p2399,p2403,p2428,p2429);
FA fa796(p2405,p2407,p2409,p2430,p2431);
FA fa797(p2415,p2417,p2419,p2432,p2433);
FA fa798(p2276,p2282,p2284,p2434,p2435);
FA fa799(p2300,p2302,p2411,p2436,p2437);
FA fa800(p2413,p2423,p2425,p2438,p2439);
HA ha419(p2290,p2292,p2440,p2441);
HA ha420(p2294,p2310,p2442,p2443);
FA fa801(p2316,p2421,p2427,p2444,p2445);
HA ha421(p2429,p2431,p2446,p2447);
FA fa802(p2433,p2304,p2306,p2448,p2449);
HA ha422(p2308,p2322,p2450,p2451);
HA ha423(p2435,p2437,p2452,p2453);
FA fa803(p2439,p2441,p2443,p2454,p2455);
HA ha424(p2447,p2312,p2456,p2457);
FA fa804(p2314,p2318,p2445,p2458,p2459);
FA fa805(p2451,p2453,p2320,p2460,p2461);
HA ha425(p2324,p2449,p2462,p2463);
FA fa806(p2455,p2457,p2326,p2464,p2465);
HA ha426(p2328,p2330,p2466,p2467);
FA fa807(p2459,p2461,p2463,p2468,p2469);
FA fa808(p2332,p2334,p2465,p2470,p2471);
FA fa809(p2467,p2336,p2338,p2472,p2473);
HA ha427(p2469,p2340,p2474,p2475);
FA fa810(p2342,p2471,p2344,p2476,p2477);
FA fa811(p2350,p2473,p2475,p2478,p2479);
HA ha428(p2346,p2352,p2480,p2481);
FA fa812(p2354,p2477,p2348,p2482,p2483);
FA fa813(p2479,p2481,p2483,p2484,p2485);
HA ha429(p2356,p2485,p2486,p2487);
HA ha430(p2358,p2360,p2488,p2489);
FA fa814(p2487,p2489,p2362,p2490,p2491);
FA fa815(ip_0_43,ip_1_42,ip_2_41,p2492,p2493);
FA fa816(ip_3_40,ip_4_39,ip_5_38,p2494,p2495);
FA fa817(ip_6_37,ip_7_36,ip_8_35,p2496,p2497);
HA ha431(ip_9_34,ip_10_33,p2498,p2499);
FA fa818(ip_11_32,ip_12_31,ip_13_30,p2500,p2501);
HA ha432(ip_14_29,ip_15_28,p2502,p2503);
FA fa819(ip_16_27,ip_17_26,ip_18_25,p2504,p2505);
FA fa820(ip_19_24,ip_20_23,ip_21_22,p2506,p2507);
FA fa821(ip_22_21,ip_23_20,ip_24_19,p2508,p2509);
HA ha433(ip_25_18,ip_26_17,p2510,p2511);
FA fa822(ip_27_16,ip_28_15,ip_29_14,p2512,p2513);
HA ha434(ip_30_13,ip_31_12,p2514,p2515);
FA fa823(ip_32_11,ip_33_10,ip_34_9,p2516,p2517);
FA fa824(ip_35_8,ip_36_7,ip_37_6,p2518,p2519);
FA fa825(ip_38_5,ip_39_4,ip_40_3,p2520,p2521);
HA ha435(ip_41_2,ip_42_1,p2522,p2523);
FA fa826(ip_43_0,p2364,p2366,p2524,p2525);
FA fa827(p2370,p2382,p2390,p2526,p2527);
FA fa828(p2499,p2503,p2511,p2528,p2529);
HA ha436(p2515,p2523,p2530,p2531);
HA ha437(p2400,p2493,p2532,p2533);
FA fa829(p2495,p2497,p2501,p2534,p2535);
FA fa830(p2505,p2507,p2509,p2536,p2537);
HA ha438(p2513,p2517,p2538,p2539);
FA fa831(p2519,p2521,p2531,p2540,p2541);
FA fa832(p2368,p2372,p2374,p2542,p2543);
FA fa833(p2376,p2378,p2380,p2544,p2545);
FA fa834(p2384,p2386,p2388,p2546,p2547);
FA fa835(p2392,p2394,p2406,p2548,p2549);
FA fa836(p2408,p2414,p2416,p2550,p2551);
FA fa837(p2418,p2525,p2527,p2552,p2553);
FA fa838(p2529,p2533,p2539,p2554,p2555);
FA fa839(p2396,p2398,p2402,p2556,p2557);
FA fa840(p2404,p2422,p2424,p2558,p2559);
FA fa841(p2535,p2537,p2541,p2560,p2561);
FA fa842(p2410,p2412,p2543,p2562,p2563);
FA fa843(p2545,p2547,p2549,p2564,p2565);
HA ha439(p2551,p2553,p2566,p2567);
FA fa844(p2555,p2420,p2426,p2568,p2569);
HA ha440(p2428,p2430,p2570,p2571);
FA fa845(p2432,p2440,p2442,p2572,p2573);
FA fa846(p2446,p2557,p2559,p2574,p2575);
HA ha441(p2561,p2567,p2576,p2577);
FA fa847(p2434,p2436,p2438,p2578,p2579);
FA fa848(p2450,p2452,p2563,p2580,p2581);
HA ha442(p2565,p2571,p2582,p2583);
HA ha443(p2577,p2444,p2584,p2585);
HA ha444(p2456,p2569,p2586,p2587);
HA ha445(p2573,p2575,p2588,p2589);
FA fa849(p2583,p2448,p2454,p2590,p2591);
HA ha446(p2462,p2579,p2592,p2593);
HA ha447(p2581,p2585,p2594,p2595);
FA fa850(p2587,p2589,p2458,p2596,p2597);
HA ha448(p2460,p2466,p2598,p2599);
HA ha449(p2593,p2595,p2600,p2601);
FA fa851(p2464,p2591,p2597,p2602,p2603);
FA fa852(p2599,p2601,p2468,p2604,p2605);
FA fa853(p2470,p2474,p2603,p2606,p2607);
HA ha450(p2605,p2472,p2608,p2609);
HA ha451(p2476,p2480,p2610,p2611);
FA fa854(p2607,p2609,p2478,p2612,p2613);
FA fa855(p2611,p2482,p2613,p2614,p2615);
HA ha452(p2484,p2486,p2616,p2617);
FA fa856(p2488,p2615,p2617,p2618,p2619);
HA ha453(ip_0_44,ip_1_43,p2620,p2621);
FA fa857(ip_2_42,ip_3_41,ip_4_40,p2622,p2623);
FA fa858(ip_5_39,ip_6_38,ip_7_37,p2624,p2625);
FA fa859(ip_8_36,ip_9_35,ip_10_34,p2626,p2627);
FA fa860(ip_11_33,ip_12_32,ip_13_31,p2628,p2629);
FA fa861(ip_14_30,ip_15_29,ip_16_28,p2630,p2631);
FA fa862(ip_17_27,ip_18_26,ip_19_25,p2632,p2633);
FA fa863(ip_20_24,ip_21_23,ip_22_22,p2634,p2635);
FA fa864(ip_23_21,ip_24_20,ip_25_19,p2636,p2637);
HA ha454(ip_26_18,ip_27_17,p2638,p2639);
FA fa865(ip_28_16,ip_29_15,ip_30_14,p2640,p2641);
HA ha455(ip_31_13,ip_32_12,p2642,p2643);
HA ha456(ip_33_11,ip_34_10,p2644,p2645);
FA fa866(ip_35_9,ip_36_8,ip_37_7,p2646,p2647);
FA fa867(ip_38_6,ip_39_5,ip_40_4,p2648,p2649);
HA ha457(ip_41_3,ip_42_2,p2650,p2651);
HA ha458(ip_43_1,ip_44_0,p2652,p2653);
FA fa868(p2498,p2502,p2510,p2654,p2655);
HA ha459(p2514,p2522,p2656,p2657);
FA fa869(p2621,p2639,p2643,p2658,p2659);
FA fa870(p2645,p2651,p2653,p2660,p2661);
HA ha460(p2530,p2623,p2662,p2663);
FA fa871(p2625,p2627,p2629,p2664,p2665);
FA fa872(p2631,p2633,p2635,p2666,p2667);
FA fa873(p2637,p2641,p2647,p2668,p2669);
FA fa874(p2649,p2657,p2492,p2670,p2671);
FA fa875(p2494,p2496,p2500,p2672,p2673);
FA fa876(p2504,p2506,p2508,p2674,p2675);
FA fa877(p2512,p2516,p2518,p2676,p2677);
HA ha461(p2520,p2532,p2678,p2679);
HA ha462(p2538,p2655,p2680,p2681);
HA ha463(p2659,p2661,p2682,p2683);
FA fa878(p2663,p2524,p2526,p2684,p2685);
FA fa879(p2528,p2665,p2667,p2686,p2687);
FA fa880(p2669,p2671,p2679,p2688,p2689);
FA fa881(p2681,p2683,p2534,p2690,p2691);
FA fa882(p2536,p2540,p2673,p2692,p2693);
HA ha464(p2675,p2677,p2694,p2695);
HA ha465(p2542,p2544,p2696,p2697);
HA ha466(p2546,p2548,p2698,p2699);
FA fa883(p2550,p2552,p2554,p2700,p2701);
HA ha467(p2566,p2685,p2702,p2703);
HA ha468(p2687,p2689,p2704,p2705);
HA ha469(p2691,p2695,p2706,p2707);
FA fa884(p2556,p2558,p2560,p2708,p2709);
HA ha470(p2570,p2576,p2710,p2711);
FA fa885(p2693,p2697,p2699,p2712,p2713);
FA fa886(p2703,p2705,p2707,p2714,p2715);
FA fa887(p2562,p2564,p2582,p2716,p2717);
HA ha471(p2701,p2711,p2718,p2719);
HA ha472(p2568,p2572,p2720,p2721);
FA fa888(p2574,p2584,p2586,p2722,p2723);
FA fa889(p2588,p2709,p2713,p2724,p2725);
HA ha473(p2715,p2719,p2726,p2727);
FA fa890(p2578,p2580,p2592,p2728,p2729);
HA ha474(p2594,p2717,p2730,p2731);
HA ha475(p2721,p2727,p2732,p2733);
FA fa891(p2598,p2600,p2723,p2734,p2735);
FA fa892(p2725,p2731,p2733,p2736,p2737);
HA ha476(p2590,p2596,p2738,p2739);
FA fa893(p2729,p2735,p2737,p2740,p2741);
HA ha477(p2739,p2602,p2742,p2743);
FA fa894(p2604,p2608,p2741,p2744,p2745);
FA fa895(p2743,p2606,p2610,p2746,p2747);
HA ha478(p2745,p2612,p2748,p2749);
HA ha479(p2747,p2616,p2750,p2751);
FA fa896(p2749,p2614,p2751,p2752,p2753);
HA ha480(ip_0_45,ip_1_44,p2754,p2755);
FA fa897(ip_2_43,ip_3_42,ip_4_41,p2756,p2757);
FA fa898(ip_5_40,ip_6_39,ip_7_38,p2758,p2759);
HA ha481(ip_8_37,ip_9_36,p2760,p2761);
HA ha482(ip_10_35,ip_11_34,p2762,p2763);
HA ha483(ip_12_33,ip_13_32,p2764,p2765);
HA ha484(ip_14_31,ip_15_30,p2766,p2767);
HA ha485(ip_16_29,ip_17_28,p2768,p2769);
HA ha486(ip_18_27,ip_19_26,p2770,p2771);
HA ha487(ip_20_25,ip_21_24,p2772,p2773);
HA ha488(ip_22_23,ip_23_22,p2774,p2775);
FA fa899(ip_24_21,ip_25_20,ip_26_19,p2776,p2777);
HA ha489(ip_27_18,ip_28_17,p2778,p2779);
FA fa900(ip_29_16,ip_30_15,ip_31_14,p2780,p2781);
FA fa901(ip_32_13,ip_33_12,ip_34_11,p2782,p2783);
FA fa902(ip_35_10,ip_36_9,ip_37_8,p2784,p2785);
FA fa903(ip_38_7,ip_39_6,ip_40_5,p2786,p2787);
FA fa904(ip_41_4,ip_42_3,ip_43_2,p2788,p2789);
FA fa905(ip_44_1,ip_45_0,p2620,p2790,p2791);
FA fa906(p2638,p2642,p2644,p2792,p2793);
FA fa907(p2650,p2652,p2755,p2794,p2795);
HA ha490(p2761,p2763,p2796,p2797);
FA fa908(p2765,p2767,p2769,p2798,p2799);
HA ha491(p2771,p2773,p2800,p2801);
HA ha492(p2775,p2779,p2802,p2803);
FA fa909(p2656,p2757,p2759,p2804,p2805);
FA fa910(p2777,p2781,p2783,p2806,p2807);
FA fa911(p2785,p2787,p2789,p2808,p2809);
HA ha493(p2791,p2797,p2810,p2811);
FA fa912(p2801,p2803,p2622,p2812,p2813);
HA ha494(p2624,p2626,p2814,p2815);
FA fa913(p2628,p2630,p2632,p2816,p2817);
HA ha495(p2634,p2636,p2818,p2819);
FA fa914(p2640,p2646,p2648,p2820,p2821);
HA ha496(p2662,p2793,p2822,p2823);
HA ha497(p2795,p2799,p2824,p2825);
HA ha498(p2811,p2654,p2826,p2827);
HA ha499(p2658,p2660,p2828,p2829);
FA fa915(p2678,p2680,p2682,p2830,p2831);
FA fa916(p2805,p2807,p2809,p2832,p2833);
HA ha500(p2813,p2815,p2834,p2835);
FA fa917(p2819,p2823,p2825,p2836,p2837);
HA ha501(p2664,p2666,p2838,p2839);
FA fa918(p2668,p2670,p2817,p2840,p2841);
FA fa919(p2821,p2827,p2829,p2842,p2843);
FA fa920(p2835,p2672,p2674,p2844,p2845);
FA fa921(p2676,p2694,p2831,p2846,p2847);
FA fa922(p2833,p2837,p2839,p2848,p2849);
FA fa923(p2684,p2686,p2688,p2850,p2851);
HA ha502(p2690,p2696,p2852,p2853);
FA fa924(p2698,p2702,p2704,p2854,p2855);
FA fa925(p2706,p2841,p2843,p2856,p2857);
HA ha503(p2692,p2710,p2858,p2859);
FA fa926(p2845,p2847,p2849,p2860,p2861);
FA fa927(p2853,p2700,p2718,p2862,p2863);
FA fa928(p2851,p2855,p2857,p2864,p2865);
HA ha504(p2859,p2708,p2866,p2867);
FA fa929(p2712,p2714,p2720,p2868,p2869);
FA fa930(p2726,p2861,p2716,p2870,p2871);
HA ha505(p2730,p2732,p2872,p2873);
HA ha506(p2863,p2865,p2874,p2875);
FA fa931(p2867,p2722,p2724,p2876,p2877);
HA ha507(p2869,p2871,p2878,p2879);
FA fa932(p2873,p2875,p2728,p2880,p2881);
HA ha508(p2738,p2879,p2882,p2883);
HA ha509(p2734,p2736,p2884,p2885);
FA fa933(p2877,p2881,p2883,p2886,p2887);
HA ha510(p2742,p2885,p2888,p2889);
HA ha511(p2740,p2887,p2890,p2891);
FA fa934(p2889,p2891,p2744,p2892,p2893);
FA fa935(p2746,p2748,p2893,p2894,p2895);
FA fa936(p2750,p2895,p2752,p2896,p2897);
HA ha512(ip_0_46,ip_1_45,p2898,p2899);
FA fa937(ip_2_44,ip_3_43,ip_4_42,p2900,p2901);
FA fa938(ip_5_41,ip_6_40,ip_7_39,p2902,p2903);
HA ha513(ip_8_38,ip_9_37,p2904,p2905);
FA fa939(ip_10_36,ip_11_35,ip_12_34,p2906,p2907);
FA fa940(ip_13_33,ip_14_32,ip_15_31,p2908,p2909);
HA ha514(ip_16_30,ip_17_29,p2910,p2911);
FA fa941(ip_18_28,ip_19_27,ip_20_26,p2912,p2913);
FA fa942(ip_21_25,ip_22_24,ip_23_23,p2914,p2915);
HA ha515(ip_24_22,ip_25_21,p2916,p2917);
HA ha516(ip_26_20,ip_27_19,p2918,p2919);
FA fa943(ip_28_18,ip_29_17,ip_30_16,p2920,p2921);
FA fa944(ip_31_15,ip_32_14,ip_33_13,p2922,p2923);
FA fa945(ip_34_12,ip_35_11,ip_36_10,p2924,p2925);
FA fa946(ip_37_9,ip_38_8,ip_39_7,p2926,p2927);
FA fa947(ip_40_6,ip_41_5,ip_42_4,p2928,p2929);
FA fa948(ip_43_3,ip_44_2,ip_45_1,p2930,p2931);
FA fa949(ip_46_0,p2754,p2760,p2932,p2933);
FA fa950(p2762,p2764,p2766,p2934,p2935);
HA ha517(p2768,p2770,p2936,p2937);
HA ha518(p2772,p2774,p2938,p2939);
HA ha519(p2778,p2899,p2940,p2941);
HA ha520(p2905,p2911,p2942,p2943);
HA ha521(p2917,p2919,p2944,p2945);
FA fa951(p2796,p2800,p2802,p2946,p2947);
FA fa952(p2901,p2903,p2907,p2948,p2949);
FA fa953(p2909,p2913,p2915,p2950,p2951);
FA fa954(p2921,p2923,p2925,p2952,p2953);
FA fa955(p2927,p2929,p2931,p2954,p2955);
HA ha522(p2937,p2939,p2956,p2957);
HA ha523(p2941,p2943,p2958,p2959);
FA fa956(p2945,p2756,p2758,p2960,p2961);
FA fa957(p2776,p2780,p2782,p2962,p2963);
FA fa958(p2784,p2786,p2788,p2964,p2965);
FA fa959(p2790,p2810,p2933,p2966,p2967);
HA ha524(p2935,p2957,p2968,p2969);
HA ha525(p2959,p2792,p2970,p2971);
FA fa960(p2794,p2798,p2814,p2972,p2973);
FA fa961(p2818,p2822,p2824,p2974,p2975);
FA fa962(p2947,p2949,p2951,p2976,p2977);
FA fa963(p2953,p2955,p2969,p2978,p2979);
FA fa964(p2804,p2806,p2808,p2980,p2981);
HA ha526(p2812,p2826,p2982,p2983);
HA ha527(p2828,p2834,p2984,p2985);
HA ha528(p2961,p2963,p2986,p2987);
HA ha529(p2965,p2967,p2988,p2989);
FA fa965(p2971,p2816,p2820,p2990,p2991);
FA fa966(p2838,p2973,p2975,p2992,p2993);
FA fa967(p2977,p2979,p2983,p2994,p2995);
FA fa968(p2985,p2987,p2989,p2996,p2997);
FA fa969(p2830,p2832,p2836,p2998,p2999);
FA fa970(p2981,p2840,p2842,p3000,p3001);
FA fa971(p2852,p2991,p2993,p3002,p3003);
HA ha530(p2995,p2997,p3004,p3005);
FA fa972(p2844,p2846,p2848,p3006,p3007);
FA fa973(p2858,p2999,p3005,p3008,p3009);
HA ha531(p2850,p2854,p3010,p3011);
FA fa974(p2856,p3001,p3003,p3012,p3013);
FA fa975(p2860,p2866,p3007,p3014,p3015);
FA fa976(p3009,p3011,p2862,p3016,p3017);
FA fa977(p2864,p2872,p2874,p3018,p3019);
FA fa978(p3013,p2868,p2870,p3020,p3021);
FA fa979(p2878,p3015,p3017,p3022,p3023);
HA ha532(p2882,p3019,p3024,p3025);
HA ha533(p2876,p2880,p3026,p3027);
FA fa980(p2884,p3021,p3023,p3028,p3029);
HA ha534(p3025,p2888,p3030,p3031);
FA fa981(p3027,p2886,p2890,p3032,p3033);
FA fa982(p3029,p3031,p3033,p3034,p3035);
FA fa983(p2892,p3035,p2894,p3036,p3037);
FA fa984(ip_0_47,ip_1_46,ip_2_45,p3038,p3039);
FA fa985(ip_3_44,ip_4_43,ip_5_42,p3040,p3041);
HA ha535(ip_6_41,ip_7_40,p3042,p3043);
HA ha536(ip_8_39,ip_9_38,p3044,p3045);
FA fa986(ip_10_37,ip_11_36,ip_12_35,p3046,p3047);
FA fa987(ip_13_34,ip_14_33,ip_15_32,p3048,p3049);
FA fa988(ip_16_31,ip_17_30,ip_18_29,p3050,p3051);
HA ha537(ip_19_28,ip_20_27,p3052,p3053);
FA fa989(ip_21_26,ip_22_25,ip_23_24,p3054,p3055);
FA fa990(ip_24_23,ip_25_22,ip_26_21,p3056,p3057);
FA fa991(ip_27_20,ip_28_19,ip_29_18,p3058,p3059);
FA fa992(ip_30_17,ip_31_16,ip_32_15,p3060,p3061);
FA fa993(ip_33_14,ip_34_13,ip_35_12,p3062,p3063);
HA ha538(ip_36_11,ip_37_10,p3064,p3065);
FA fa994(ip_38_9,ip_39_8,ip_40_7,p3066,p3067);
HA ha539(ip_41_6,ip_42_5,p3068,p3069);
HA ha540(ip_43_4,ip_44_3,p3070,p3071);
FA fa995(ip_45_2,ip_46_1,ip_47_0,p3072,p3073);
FA fa996(p2898,p2904,p2910,p3074,p3075);
HA ha541(p2916,p2918,p3076,p3077);
FA fa997(p3043,p3045,p3053,p3078,p3079);
HA ha542(p3065,p3069,p3080,p3081);
HA ha543(p3071,p2936,p3082,p3083);
FA fa998(p2938,p2940,p2942,p3084,p3085);
FA fa999(p2944,p3039,p3041,p3086,p3087);
HA ha544(p3047,p3049,p3088,p3089);
FA fa1000(p3051,p3055,p3057,p3090,p3091);
FA fa1001(p3059,p3061,p3063,p3092,p3093);
FA fa1002(p3067,p3073,p3077,p3094,p3095);
FA fa1003(p3081,p2900,p2902,p3096,p3097);
FA fa1004(p2906,p2908,p2912,p3098,p3099);
FA fa1005(p2914,p2920,p2922,p3100,p3101);
FA fa1006(p2924,p2926,p2928,p3102,p3103);
FA fa1007(p2930,p2956,p2958,p3104,p3105);
HA ha545(p3075,p3079,p3106,p3107);
HA ha546(p3083,p3089,p3108,p3109);
FA fa1008(p2932,p2934,p2968,p3110,p3111);
FA fa1009(p3085,p3087,p3091,p3112,p3113);
HA ha547(p3093,p3095,p3114,p3115);
FA fa1010(p3107,p3109,p2946,p3116,p3117);
FA fa1011(p2948,p2950,p2952,p3118,p3119);
FA fa1012(p2954,p2970,p3097,p3120,p3121);
HA ha548(p3099,p3101,p3122,p3123);
HA ha549(p3103,p3105,p3124,p3125);
HA ha550(p3115,p2960,p3126,p3127);
FA fa1013(p2962,p2964,p2966,p3128,p3129);
FA fa1014(p2982,p2984,p2986,p3130,p3131);
FA fa1015(p2988,p3111,p3113,p3132,p3133);
HA ha551(p3117,p3123,p3134,p3135);
FA fa1016(p3125,p2972,p2974,p3136,p3137);
HA ha552(p2976,p2978,p3138,p3139);
FA fa1017(p3119,p3121,p3127,p3140,p3141);
HA ha553(p3135,p2980,p3142,p3143);
FA fa1018(p3129,p3131,p3133,p3144,p3145);
FA fa1019(p3139,p2990,p2992,p3146,p3147);
HA ha554(p2994,p2996,p3148,p3149);
FA fa1020(p3004,p3137,p3141,p3150,p3151);
FA fa1021(p3143,p2998,p3145,p3152,p3153);
FA fa1022(p3149,p3000,p3002,p3154,p3155);
FA fa1023(p3010,p3147,p3151,p3156,p3157);
FA fa1024(p3006,p3008,p3153,p3158,p3159);
FA fa1025(p3012,p3155,p3157,p3160,p3161);
FA fa1026(p3014,p3016,p3159,p3162,p3163);
FA fa1027(p3018,p3024,p3161,p3164,p3165);
FA fa1028(p3020,p3022,p3026,p3166,p3167);
FA fa1029(p3163,p3030,p3165,p3168,p3169);
FA fa1030(p3028,p3167,p3169,p3170,p3171);
HA ha555(p3032,p3171,p3172,p3173);
FA fa1031(p3034,p3173,p3036,p3174,p3175);
FA fa1032(ip_0_48,ip_1_47,ip_2_46,p3176,p3177);
FA fa1033(ip_3_45,ip_4_44,ip_5_43,p3178,p3179);
FA fa1034(ip_6_42,ip_7_41,ip_8_40,p3180,p3181);
HA ha556(ip_9_39,ip_10_38,p3182,p3183);
FA fa1035(ip_11_37,ip_12_36,ip_13_35,p3184,p3185);
FA fa1036(ip_14_34,ip_15_33,ip_16_32,p3186,p3187);
FA fa1037(ip_17_31,ip_18_30,ip_19_29,p3188,p3189);
FA fa1038(ip_20_28,ip_21_27,ip_22_26,p3190,p3191);
HA ha557(ip_23_25,ip_24_24,p3192,p3193);
HA ha558(ip_25_23,ip_26_22,p3194,p3195);
HA ha559(ip_27_21,ip_28_20,p3196,p3197);
HA ha560(ip_29_19,ip_30_18,p3198,p3199);
FA fa1039(ip_31_17,ip_32_16,ip_33_15,p3200,p3201);
FA fa1040(ip_34_14,ip_35_13,ip_36_12,p3202,p3203);
HA ha561(ip_37_11,ip_38_10,p3204,p3205);
FA fa1041(ip_39_9,ip_40_8,ip_41_7,p3206,p3207);
FA fa1042(ip_42_6,ip_43_5,ip_44_4,p3208,p3209);
FA fa1043(ip_45_3,ip_46_2,ip_47_1,p3210,p3211);
FA fa1044(ip_48_0,p3042,p3044,p3212,p3213);
FA fa1045(p3052,p3064,p3068,p3214,p3215);
HA ha562(p3070,p3183,p3216,p3217);
HA ha563(p3193,p3195,p3218,p3219);
HA ha564(p3197,p3199,p3220,p3221);
FA fa1046(p3205,p3076,p3080,p3222,p3223);
HA ha565(p3177,p3179,p3224,p3225);
FA fa1047(p3181,p3185,p3187,p3226,p3227);
HA ha566(p3189,p3191,p3228,p3229);
FA fa1048(p3201,p3203,p3207,p3230,p3231);
FA fa1049(p3209,p3211,p3217,p3232,p3233);
HA ha567(p3219,p3221,p3234,p3235);
HA ha568(p3038,p3040,p3236,p3237);
FA fa1050(p3046,p3048,p3050,p3238,p3239);
FA fa1051(p3054,p3056,p3058,p3240,p3241);
HA ha569(p3060,p3062,p3242,p3243);
HA ha570(p3066,p3072,p3244,p3245);
HA ha571(p3082,p3088,p3246,p3247);
FA fa1052(p3213,p3215,p3225,p3248,p3249);
FA fa1053(p3229,p3235,p3074,p3250,p3251);
HA ha572(p3078,p3106,p3252,p3253);
FA fa1054(p3108,p3223,p3227,p3254,p3255);
FA fa1055(p3231,p3233,p3237,p3256,p3257);
FA fa1056(p3243,p3245,p3247,p3258,p3259);
FA fa1057(p3084,p3086,p3090,p3260,p3261);
HA ha573(p3092,p3094,p3262,p3263);
HA ha574(p3114,p3239,p3264,p3265);
FA fa1058(p3241,p3249,p3251,p3266,p3267);
FA fa1059(p3253,p3096,p3098,p3268,p3269);
FA fa1060(p3100,p3102,p3104,p3270,p3271);
FA fa1061(p3122,p3124,p3255,p3272,p3273);
FA fa1062(p3257,p3259,p3263,p3274,p3275);
FA fa1063(p3265,p3110,p3112,p3276,p3277);
FA fa1064(p3116,p3126,p3134,p3278,p3279);
FA fa1065(p3261,p3267,p3118,p3280,p3281);
HA ha575(p3120,p3138,p3282,p3283);
FA fa1066(p3269,p3271,p3273,p3284,p3285);
HA ha576(p3275,p3128,p3286,p3287);
HA ha577(p3130,p3132,p3288,p3289);
HA ha578(p3142,p3277,p3290,p3291);
HA ha579(p3279,p3281,p3292,p3293);
HA ha580(p3283,p3136,p3294,p3295);
FA fa1067(p3140,p3148,p3285,p3296,p3297);
FA fa1068(p3287,p3289,p3291,p3298,p3299);
FA fa1069(p3293,p3144,p3295,p3300,p3301);
FA fa1070(p3146,p3150,p3297,p3302,p3303);
FA fa1071(p3299,p3152,p3301,p3304,p3305);
HA ha581(p3154,p3156,p3306,p3307);
HA ha582(p3303,p3158,p3308,p3309);
FA fa1072(p3305,p3307,p3160,p3310,p3311);
HA ha583(p3309,p3162,p3312,p3313);
HA ha584(p3311,p3164,p3314,p3315);
HA ha585(p3313,p3166,p3316,p3317);
HA ha586(p3315,p3168,p3318,p3319);
HA ha587(p3317,p3170,p3320,p3321);
FA fa1073(p3172,p3319,p3321,p3322,p3323);
HA ha588(ip_0_49,ip_1_48,p3324,p3325);
FA fa1074(ip_2_47,ip_3_46,ip_4_45,p3326,p3327);
HA ha589(ip_5_44,ip_6_43,p3328,p3329);
HA ha590(ip_7_42,ip_8_41,p3330,p3331);
HA ha591(ip_9_40,ip_10_39,p3332,p3333);
FA fa1075(ip_11_38,ip_12_37,ip_13_36,p3334,p3335);
FA fa1076(ip_14_35,ip_15_34,ip_16_33,p3336,p3337);
FA fa1077(ip_17_32,ip_18_31,ip_19_30,p3338,p3339);
FA fa1078(ip_20_29,ip_21_28,ip_22_27,p3340,p3341);
HA ha592(ip_23_26,ip_24_25,p3342,p3343);
FA fa1079(ip_25_24,ip_26_23,ip_27_22,p3344,p3345);
FA fa1080(ip_28_21,ip_29_20,ip_30_19,p3346,p3347);
FA fa1081(ip_31_18,ip_32_17,ip_33_16,p3348,p3349);
FA fa1082(ip_34_15,ip_35_14,ip_36_13,p3350,p3351);
FA fa1083(ip_37_12,ip_38_11,ip_39_10,p3352,p3353);
FA fa1084(ip_40_9,ip_41_8,ip_42_7,p3354,p3355);
HA ha593(ip_43_6,ip_44_5,p3356,p3357);
HA ha594(ip_45_4,ip_46_3,p3358,p3359);
FA fa1085(ip_47_2,ip_48_1,ip_49_0,p3360,p3361);
HA ha595(p3182,p3192,p3362,p3363);
FA fa1086(p3194,p3196,p3198,p3364,p3365);
HA ha596(p3204,p3325,p3366,p3367);
HA ha597(p3329,p3331,p3368,p3369);
HA ha598(p3333,p3343,p3370,p3371);
FA fa1087(p3357,p3359,p3216,p3372,p3373);
HA ha599(p3218,p3220,p3374,p3375);
FA fa1088(p3327,p3335,p3337,p3376,p3377);
FA fa1089(p3339,p3341,p3345,p3378,p3379);
HA ha600(p3347,p3349,p3380,p3381);
HA ha601(p3351,p3353,p3382,p3383);
FA fa1090(p3355,p3361,p3363,p3384,p3385);
FA fa1091(p3367,p3369,p3371,p3386,p3387);
FA fa1092(p3176,p3178,p3180,p3388,p3389);
FA fa1093(p3184,p3186,p3188,p3390,p3391);
FA fa1094(p3190,p3200,p3202,p3392,p3393);
HA ha602(p3206,p3208,p3394,p3395);
FA fa1095(p3210,p3224,p3228,p3396,p3397);
FA fa1096(p3234,p3365,p3373,p3398,p3399);
HA ha603(p3375,p3381,p3400,p3401);
FA fa1097(p3383,p3212,p3214,p3402,p3403);
FA fa1098(p3236,p3242,p3244,p3404,p3405);
FA fa1099(p3246,p3377,p3379,p3406,p3407);
FA fa1100(p3385,p3387,p3395,p3408,p3409);
FA fa1101(p3401,p3222,p3226,p3410,p3411);
HA ha604(p3230,p3232,p3412,p3413);
FA fa1102(p3252,p3389,p3391,p3414,p3415);
FA fa1103(p3393,p3397,p3399,p3416,p3417);
FA fa1104(p3238,p3240,p3248,p3418,p3419);
FA fa1105(p3250,p3262,p3264,p3420,p3421);
FA fa1106(p3403,p3405,p3407,p3422,p3423);
HA ha605(p3409,p3413,p3424,p3425);
HA ha606(p3254,p3256,p3426,p3427);
FA fa1107(p3258,p3411,p3415,p3428,p3429);
FA fa1108(p3417,p3425,p3260,p3430,p3431);
HA ha607(p3266,p3419,p3432,p3433);
FA fa1109(p3421,p3423,p3427,p3434,p3435);
HA ha608(p3268,p3270,p3436,p3437);
HA ha609(p3272,p3274,p3438,p3439);
FA fa1110(p3282,p3429,p3431,p3440,p3441);
HA ha610(p3433,p3276,p3442,p3443);
FA fa1111(p3278,p3280,p3286,p3444,p3445);
HA ha611(p3288,p3290,p3446,p3447);
FA fa1112(p3292,p3435,p3437,p3448,p3449);
FA fa1113(p3439,p3284,p3294,p3450,p3451);
FA fa1114(p3441,p3443,p3447,p3452,p3453);
FA fa1115(p3445,p3449,p3296,p3454,p3455);
FA fa1116(p3298,p3451,p3453,p3456,p3457);
FA fa1117(p3300,p3455,p3302,p3458,p3459);
HA ha612(p3306,p3457,p3460,p3461);
FA fa1118(p3304,p3308,p3459,p3462,p3463);
FA fa1119(p3461,p3310,p3312,p3464,p3465);
HA ha613(p3463,p3314,p3466,p3467);
FA fa1120(p3316,p3465,p3467,p3468,p3469);
HA ha614(p3318,p3320,p3470,p3471);
HA ha615(p3469,p3471,p3472,p3473);
FA fa1121(ip_0_50,ip_1_49,ip_2_48,p3474,p3475);
FA fa1122(ip_3_47,ip_4_46,ip_5_45,p3476,p3477);
FA fa1123(ip_6_44,ip_7_43,ip_8_42,p3478,p3479);
FA fa1124(ip_9_41,ip_10_40,ip_11_39,p3480,p3481);
FA fa1125(ip_12_38,ip_13_37,ip_14_36,p3482,p3483);
FA fa1126(ip_15_35,ip_16_34,ip_17_33,p3484,p3485);
HA ha616(ip_18_32,ip_19_31,p3486,p3487);
FA fa1127(ip_20_30,ip_21_29,ip_22_28,p3488,p3489);
HA ha617(ip_23_27,ip_24_26,p3490,p3491);
FA fa1128(ip_25_25,ip_26_24,ip_27_23,p3492,p3493);
HA ha618(ip_28_22,ip_29_21,p3494,p3495);
HA ha619(ip_30_20,ip_31_19,p3496,p3497);
FA fa1129(ip_32_18,ip_33_17,ip_34_16,p3498,p3499);
HA ha620(ip_35_15,ip_36_14,p3500,p3501);
HA ha621(ip_37_13,ip_38_12,p3502,p3503);
FA fa1130(ip_39_11,ip_40_10,ip_41_9,p3504,p3505);
FA fa1131(ip_42_8,ip_43_7,ip_44_6,p3506,p3507);
HA ha622(ip_45_5,ip_46_4,p3508,p3509);
HA ha623(ip_47_3,ip_48_2,p3510,p3511);
HA ha624(ip_49_1,ip_50_0,p3512,p3513);
FA fa1132(p3324,p3328,p3330,p3514,p3515);
FA fa1133(p3332,p3342,p3356,p3516,p3517);
HA ha625(p3358,p3487,p3518,p3519);
HA ha626(p3491,p3495,p3520,p3521);
FA fa1134(p3497,p3501,p3503,p3522,p3523);
FA fa1135(p3509,p3511,p3513,p3524,p3525);
FA fa1136(p3362,p3366,p3368,p3526,p3527);
HA ha627(p3370,p3475,p3528,p3529);
HA ha628(p3477,p3479,p3530,p3531);
FA fa1137(p3481,p3483,p3485,p3532,p3533);
HA ha629(p3489,p3493,p3534,p3535);
FA fa1138(p3499,p3505,p3507,p3536,p3537);
FA fa1139(p3519,p3521,p3326,p3538,p3539);
FA fa1140(p3334,p3336,p3338,p3540,p3541);
FA fa1141(p3340,p3344,p3346,p3542,p3543);
FA fa1142(p3348,p3350,p3352,p3544,p3545);
HA ha630(p3354,p3360,p3546,p3547);
FA fa1143(p3374,p3380,p3382,p3548,p3549);
FA fa1144(p3515,p3517,p3523,p3550,p3551);
FA fa1145(p3525,p3529,p3531,p3552,p3553);
FA fa1146(p3535,p3364,p3372,p3554,p3555);
FA fa1147(p3394,p3400,p3527,p3556,p3557);
HA ha631(p3533,p3537,p3558,p3559);
FA fa1148(p3539,p3547,p3376,p3560,p3561);
FA fa1149(p3378,p3384,p3386,p3562,p3563);
FA fa1150(p3541,p3543,p3545,p3564,p3565);
FA fa1151(p3549,p3551,p3553,p3566,p3567);
FA fa1152(p3559,p3388,p3390,p3568,p3569);
HA ha632(p3392,p3396,p3570,p3571);
HA ha633(p3398,p3412,p3572,p3573);
HA ha634(p3555,p3557,p3574,p3575);
HA ha635(p3561,p3402,p3576,p3577);
FA fa1153(p3404,p3406,p3408,p3578,p3579);
FA fa1154(p3424,p3563,p3565,p3580,p3581);
FA fa1155(p3567,p3571,p3573,p3582,p3583);
FA fa1156(p3575,p3410,p3414,p3584,p3585);
FA fa1157(p3416,p3426,p3569,p3586,p3587);
HA ha636(p3577,p3418,p3588,p3589);
HA ha637(p3420,p3422,p3590,p3591);
HA ha638(p3432,p3579,p3592,p3593);
FA fa1158(p3581,p3583,p3428,p3594,p3595);
FA fa1159(p3430,p3436,p3438,p3596,p3597);
FA fa1160(p3585,p3587,p3589,p3598,p3599);
FA fa1161(p3591,p3593,p3434,p3600,p3601);
FA fa1162(p3442,p3446,p3595,p3602,p3603);
FA fa1163(p3440,p3597,p3599,p3604,p3605);
HA ha639(p3601,p3444,p3606,p3607);
FA fa1164(p3448,p3603,p3450,p3608,p3609);
FA fa1165(p3452,p3605,p3607,p3610,p3611);
FA fa1166(p3454,p3609,p3456,p3612,p3613);
FA fa1167(p3460,p3611,p3458,p3614,p3615);
FA fa1168(p3613,p3615,p3462,p3616,p3617);
HA ha640(p3466,p3617,p3618,p3619);
HA ha641(p3464,p3619,p3620,p3621);
FA fa1169(p3621,p3468,p3470,p3622,p3623);
HA ha642(ip_0_51,ip_1_50,p3624,p3625);
HA ha643(ip_2_49,ip_3_48,p3626,p3627);
FA fa1170(ip_4_47,ip_5_46,ip_6_45,p3628,p3629);
HA ha644(ip_7_44,ip_8_43,p3630,p3631);
FA fa1171(ip_9_42,ip_10_41,ip_11_40,p3632,p3633);
HA ha645(ip_12_39,ip_13_38,p3634,p3635);
FA fa1172(ip_14_37,ip_15_36,ip_16_35,p3636,p3637);
FA fa1173(ip_17_34,ip_18_33,ip_19_32,p3638,p3639);
FA fa1174(ip_20_31,ip_21_30,ip_22_29,p3640,p3641);
FA fa1175(ip_23_28,ip_24_27,ip_25_26,p3642,p3643);
FA fa1176(ip_26_25,ip_27_24,ip_28_23,p3644,p3645);
HA ha646(ip_29_22,ip_30_21,p3646,p3647);
HA ha647(ip_31_20,ip_32_19,p3648,p3649);
FA fa1177(ip_33_18,ip_34_17,ip_35_16,p3650,p3651);
FA fa1178(ip_36_15,ip_37_14,ip_38_13,p3652,p3653);
HA ha648(ip_39_12,ip_40_11,p3654,p3655);
FA fa1179(ip_41_10,ip_42_9,ip_43_8,p3656,p3657);
HA ha649(ip_44_7,ip_45_6,p3658,p3659);
FA fa1180(ip_46_5,ip_47_4,ip_48_3,p3660,p3661);
FA fa1181(ip_49_2,ip_50_1,ip_51_0,p3662,p3663);
FA fa1182(p3486,p3490,p3494,p3664,p3665);
FA fa1183(p3496,p3500,p3502,p3666,p3667);
FA fa1184(p3508,p3510,p3512,p3668,p3669);
FA fa1185(p3625,p3627,p3631,p3670,p3671);
HA ha650(p3635,p3647,p3672,p3673);
FA fa1186(p3649,p3655,p3659,p3674,p3675);
HA ha651(p3518,p3520,p3676,p3677);
FA fa1187(p3629,p3633,p3637,p3678,p3679);
HA ha652(p3639,p3641,p3680,p3681);
FA fa1188(p3643,p3645,p3651,p3682,p3683);
FA fa1189(p3653,p3657,p3661,p3684,p3685);
FA fa1190(p3663,p3673,p3474,p3686,p3687);
FA fa1191(p3476,p3478,p3480,p3688,p3689);
FA fa1192(p3482,p3484,p3488,p3690,p3691);
FA fa1193(p3492,p3498,p3504,p3692,p3693);
FA fa1194(p3506,p3528,p3530,p3694,p3695);
FA fa1195(p3534,p3665,p3667,p3696,p3697);
HA ha653(p3669,p3671,p3698,p3699);
FA fa1196(p3675,p3677,p3681,p3700,p3701);
FA fa1197(p3514,p3516,p3522,p3702,p3703);
FA fa1198(p3524,p3546,p3679,p3704,p3705);
FA fa1199(p3683,p3685,p3687,p3706,p3707);
HA ha654(p3699,p3526,p3708,p3709);
FA fa1200(p3532,p3536,p3538,p3710,p3711);
HA ha655(p3558,p3689,p3712,p3713);
HA ha656(p3691,p3693,p3714,p3715);
FA fa1201(p3695,p3697,p3701,p3716,p3717);
HA ha657(p3540,p3542,p3718,p3719);
FA fa1202(p3544,p3548,p3550,p3720,p3721);
HA ha658(p3552,p3703,p3722,p3723);
FA fa1203(p3705,p3707,p3709,p3724,p3725);
HA ha659(p3713,p3715,p3726,p3727);
FA fa1204(p3554,p3556,p3560,p3728,p3729);
HA ha660(p3570,p3572,p3730,p3731);
FA fa1205(p3574,p3711,p3717,p3732,p3733);
FA fa1206(p3719,p3723,p3727,p3734,p3735);
FA fa1207(p3562,p3564,p3566,p3736,p3737);
FA fa1208(p3576,p3721,p3725,p3738,p3739);
FA fa1209(p3731,p3568,p3729,p3740,p3741);
HA ha661(p3733,p3735,p3742,p3743);
FA fa1210(p3578,p3580,p3582,p3744,p3745);
FA fa1211(p3588,p3590,p3592,p3746,p3747);
HA ha662(p3737,p3739,p3748,p3749);
FA fa1212(p3743,p3584,p3586,p3750,p3751);
FA fa1213(p3741,p3749,p3594,p3752,p3753);
FA fa1214(p3745,p3747,p3596,p3754,p3755);
FA fa1215(p3598,p3600,p3751,p3756,p3757);
FA fa1216(p3753,p3602,p3606,p3758,p3759);
FA fa1217(p3755,p3604,p3757,p3760,p3761);
FA fa1218(p3608,p3759,p3610,p3762,p3763);
HA ha663(p3761,p3612,p3764,p3765);
FA fa1219(p3763,p3614,p3765,p3766,p3767);
FA fa1220(p3616,p3618,p3767,p3768,p3769);
HA ha664(p3620,p3769,p3770,p3771);
FA fa1221(ip_0_52,ip_1_51,ip_2_50,p3772,p3773);
HA ha665(ip_3_49,ip_4_48,p3774,p3775);
HA ha666(ip_5_47,ip_6_46,p3776,p3777);
FA fa1222(ip_7_45,ip_8_44,ip_9_43,p3778,p3779);
FA fa1223(ip_10_42,ip_11_41,ip_12_40,p3780,p3781);
HA ha667(ip_13_39,ip_14_38,p3782,p3783);
HA ha668(ip_15_37,ip_16_36,p3784,p3785);
FA fa1224(ip_17_35,ip_18_34,ip_19_33,p3786,p3787);
FA fa1225(ip_20_32,ip_21_31,ip_22_30,p3788,p3789);
FA fa1226(ip_23_29,ip_24_28,ip_25_27,p3790,p3791);
HA ha669(ip_26_26,ip_27_25,p3792,p3793);
FA fa1227(ip_28_24,ip_29_23,ip_30_22,p3794,p3795);
FA fa1228(ip_31_21,ip_32_20,ip_33_19,p3796,p3797);
FA fa1229(ip_34_18,ip_35_17,ip_36_16,p3798,p3799);
HA ha670(ip_37_15,ip_38_14,p3800,p3801);
FA fa1230(ip_39_13,ip_40_12,ip_41_11,p3802,p3803);
FA fa1231(ip_42_10,ip_43_9,ip_44_8,p3804,p3805);
FA fa1232(ip_45_7,ip_46_6,ip_47_5,p3806,p3807);
FA fa1233(ip_48_4,ip_49_3,ip_50_2,p3808,p3809);
HA ha671(ip_51_1,ip_52_0,p3810,p3811);
FA fa1234(p3624,p3626,p3630,p3812,p3813);
FA fa1235(p3634,p3646,p3648,p3814,p3815);
FA fa1236(p3654,p3658,p3775,p3816,p3817);
FA fa1237(p3777,p3783,p3785,p3818,p3819);
FA fa1238(p3793,p3801,p3811,p3820,p3821);
FA fa1239(p3672,p3773,p3779,p3822,p3823);
FA fa1240(p3781,p3787,p3789,p3824,p3825);
FA fa1241(p3791,p3795,p3797,p3826,p3827);
HA ha672(p3799,p3803,p3828,p3829);
FA fa1242(p3805,p3807,p3809,p3830,p3831);
FA fa1243(p3628,p3632,p3636,p3832,p3833);
FA fa1244(p3638,p3640,p3642,p3834,p3835);
FA fa1245(p3644,p3650,p3652,p3836,p3837);
HA ha673(p3656,p3660,p3838,p3839);
HA ha674(p3662,p3676,p3840,p3841);
FA fa1246(p3680,p3813,p3815,p3842,p3843);
HA ha675(p3817,p3819,p3844,p3845);
FA fa1247(p3821,p3829,p3664,p3846,p3847);
FA fa1248(p3666,p3668,p3670,p3848,p3849);
HA ha676(p3674,p3698,p3850,p3851);
FA fa1249(p3823,p3825,p3827,p3852,p3853);
HA ha677(p3831,p3839,p3854,p3855);
HA ha678(p3841,p3845,p3856,p3857);
HA ha679(p3678,p3682,p3858,p3859);
FA fa1250(p3684,p3686,p3833,p3860,p3861);
FA fa1251(p3835,p3837,p3843,p3862,p3863);
HA ha680(p3847,p3851,p3864,p3865);
FA fa1252(p3855,p3857,p3688,p3866,p3867);
HA ha681(p3690,p3692,p3868,p3869);
HA ha682(p3694,p3696,p3870,p3871);
HA ha683(p3700,p3708,p3872,p3873);
FA fa1253(p3712,p3714,p3849,p3874,p3875);
HA ha684(p3853,p3859,p3876,p3877);
FA fa1254(p3865,p3702,p3704,p3878,p3879);
FA fa1255(p3706,p3718,p3722,p3880,p3881);
FA fa1256(p3726,p3861,p3863,p3882,p3883);
FA fa1257(p3867,p3869,p3871,p3884,p3885);
FA fa1258(p3873,p3877,p3710,p3886,p3887);
FA fa1259(p3716,p3730,p3875,p3888,p3889);
FA fa1260(p3720,p3724,p3879,p3890,p3891);
FA fa1261(p3881,p3883,p3885,p3892,p3893);
FA fa1262(p3887,p3728,p3732,p3894,p3895);
HA ha685(p3734,p3742,p3896,p3897);
FA fa1263(p3889,p3736,p3738,p3898,p3899);
HA ha686(p3748,p3891,p3900,p3901);
FA fa1264(p3893,p3897,p3740,p3902,p3903);
FA fa1265(p3895,p3901,p3744,p3904,p3905);
FA fa1266(p3746,p3899,p3903,p3906,p3907);
FA fa1267(p3750,p3752,p3905,p3908,p3909);
HA ha687(p3754,p3907,p3910,p3911);
FA fa1268(p3756,p3909,p3911,p3912,p3913);
FA fa1269(p3758,p3760,p3913,p3914,p3915);
FA fa1270(p3762,p3764,p3915,p3916,p3917);
FA fa1271(p3917,p3766,p3768,p3918,p3919);
FA fa1272(ip_0_53,ip_1_52,ip_2_51,p3920,p3921);
FA fa1273(ip_3_50,ip_4_49,ip_5_48,p3922,p3923);
FA fa1274(ip_6_47,ip_7_46,ip_8_45,p3924,p3925);
FA fa1275(ip_9_44,ip_10_43,ip_11_42,p3926,p3927);
FA fa1276(ip_12_41,ip_13_40,ip_14_39,p3928,p3929);
HA ha688(ip_15_38,ip_16_37,p3930,p3931);
FA fa1277(ip_17_36,ip_18_35,ip_19_34,p3932,p3933);
FA fa1278(ip_20_33,ip_21_32,ip_22_31,p3934,p3935);
FA fa1279(ip_23_30,ip_24_29,ip_25_28,p3936,p3937);
FA fa1280(ip_26_27,ip_27_26,ip_28_25,p3938,p3939);
FA fa1281(ip_29_24,ip_30_23,ip_31_22,p3940,p3941);
FA fa1282(ip_32_21,ip_33_20,ip_34_19,p3942,p3943);
HA ha689(ip_35_18,ip_36_17,p3944,p3945);
HA ha690(ip_37_16,ip_38_15,p3946,p3947);
FA fa1283(ip_39_14,ip_40_13,ip_41_12,p3948,p3949);
HA ha691(ip_42_11,ip_43_10,p3950,p3951);
FA fa1284(ip_44_9,ip_45_8,ip_46_7,p3952,p3953);
FA fa1285(ip_47_6,ip_48_5,ip_49_4,p3954,p3955);
FA fa1286(ip_50_3,ip_51_2,ip_52_1,p3956,p3957);
FA fa1287(ip_53_0,p3774,p3776,p3958,p3959);
FA fa1288(p3782,p3784,p3792,p3960,p3961);
HA ha692(p3800,p3810,p3962,p3963);
FA fa1289(p3931,p3945,p3947,p3964,p3965);
FA fa1290(p3951,p3921,p3923,p3966,p3967);
HA ha693(p3925,p3927,p3968,p3969);
FA fa1291(p3929,p3933,p3935,p3970,p3971);
HA ha694(p3937,p3939,p3972,p3973);
HA ha695(p3941,p3943,p3974,p3975);
HA ha696(p3949,p3953,p3976,p3977);
FA fa1292(p3955,p3957,p3963,p3978,p3979);
FA fa1293(p3772,p3778,p3780,p3980,p3981);
FA fa1294(p3786,p3788,p3790,p3982,p3983);
HA ha697(p3794,p3796,p3984,p3985);
FA fa1295(p3798,p3802,p3804,p3986,p3987);
HA ha698(p3806,p3808,p3988,p3989);
FA fa1296(p3828,p3959,p3961,p3990,p3991);
FA fa1297(p3965,p3969,p3973,p3992,p3993);
FA fa1298(p3975,p3977,p3812,p3994,p3995);
HA ha699(p3814,p3816,p3996,p3997);
FA fa1299(p3818,p3820,p3838,p3998,p3999);
FA fa1300(p3840,p3844,p3967,p4000,p4001);
FA fa1301(p3971,p3979,p3985,p4002,p4003);
FA fa1302(p3989,p3822,p3824,p4004,p4005);
FA fa1303(p3826,p3830,p3850,p4006,p4007);
HA ha700(p3854,p3856,p4008,p4009);
HA ha701(p3981,p3983,p4010,p4011);
FA fa1304(p3987,p3991,p3993,p4012,p4013);
FA fa1305(p3995,p3997,p3832,p4014,p4015);
FA fa1306(p3834,p3836,p3842,p4016,p4017);
FA fa1307(p3846,p3858,p3864,p4018,p4019);
FA fa1308(p3999,p4001,p4003,p4020,p4021);
FA fa1309(p4009,p4011,p3848,p4022,p4023);
FA fa1310(p3852,p3868,p3870,p4024,p4025);
FA fa1311(p3872,p3876,p4005,p4026,p4027);
FA fa1312(p4007,p4013,p4015,p4028,p4029);
FA fa1313(p3860,p3862,p3866,p4030,p4031);
HA ha702(p4017,p4019,p4032,p4033);
FA fa1314(p4021,p4023,p3874,p4034,p4035);
FA fa1315(p4025,p4027,p4029,p4036,p4037);
FA fa1316(p4033,p3878,p3880,p4038,p4039);
FA fa1317(p3882,p3884,p3886,p4040,p4041);
HA ha703(p4031,p4035,p4042,p4043);
HA ha704(p3888,p3896,p4044,p4045);
FA fa1318(p4037,p4043,p3890,p4046,p4047);
HA ha705(p3892,p3900,p4048,p4049);
FA fa1319(p4039,p4041,p4045,p4050,p4051);
FA fa1320(p3894,p4047,p4049,p4052,p4053);
HA ha706(p3898,p3902,p4054,p4055);
FA fa1321(p4051,p3904,p4053,p4056,p4057);
FA fa1322(p4055,p3906,p3910,p4058,p4059);
FA fa1323(p3908,p4057,p4059,p4060,p4061);
FA fa1324(p3912,p4061,p3914,p4062,p4063);
HA ha707(p3916,p4063,p4064,p4065);
HA ha708(ip_0_54,ip_1_53,p4066,p4067);
HA ha709(ip_2_52,ip_3_51,p4068,p4069);
FA fa1325(ip_4_50,ip_5_49,ip_6_48,p4070,p4071);
FA fa1326(ip_7_47,ip_8_46,ip_9_45,p4072,p4073);
HA ha710(ip_10_44,ip_11_43,p4074,p4075);
FA fa1327(ip_12_42,ip_13_41,ip_14_40,p4076,p4077);
HA ha711(ip_15_39,ip_16_38,p4078,p4079);
HA ha712(ip_17_37,ip_18_36,p4080,p4081);
FA fa1328(ip_19_35,ip_20_34,ip_21_33,p4082,p4083);
FA fa1329(ip_22_32,ip_23_31,ip_24_30,p4084,p4085);
FA fa1330(ip_25_29,ip_26_28,ip_27_27,p4086,p4087);
FA fa1331(ip_28_26,ip_29_25,ip_30_24,p4088,p4089);
FA fa1332(ip_31_23,ip_32_22,ip_33_21,p4090,p4091);
FA fa1333(ip_34_20,ip_35_19,ip_36_18,p4092,p4093);
HA ha713(ip_37_17,ip_38_16,p4094,p4095);
FA fa1334(ip_39_15,ip_40_14,ip_41_13,p4096,p4097);
HA ha714(ip_42_12,ip_43_11,p4098,p4099);
FA fa1335(ip_44_10,ip_45_9,ip_46_8,p4100,p4101);
FA fa1336(ip_47_7,ip_48_6,ip_49_5,p4102,p4103);
FA fa1337(ip_50_4,ip_51_3,ip_52_2,p4104,p4105);
FA fa1338(ip_53_1,ip_54_0,p3930,p4106,p4107);
HA ha715(p3944,p3946,p4108,p4109);
FA fa1339(p3950,p4067,p4069,p4110,p4111);
HA ha716(p4075,p4079,p4112,p4113);
FA fa1340(p4081,p4095,p4099,p4114,p4115);
FA fa1341(p3962,p4071,p4073,p4116,p4117);
HA ha717(p4077,p4083,p4118,p4119);
FA fa1342(p4085,p4087,p4089,p4120,p4121);
HA ha718(p4091,p4093,p4122,p4123);
FA fa1343(p4097,p4101,p4103,p4124,p4125);
FA fa1344(p4105,p4107,p4109,p4126,p4127);
HA ha719(p4113,p3920,p4128,p4129);
FA fa1345(p3922,p3924,p3926,p4130,p4131);
HA ha720(p3928,p3932,p4132,p4133);
FA fa1346(p3934,p3936,p3938,p4134,p4135);
FA fa1347(p3940,p3942,p3948,p4136,p4137);
HA ha721(p3952,p3954,p4138,p4139);
FA fa1348(p3956,p3968,p3972,p4140,p4141);
HA ha722(p3974,p3976,p4142,p4143);
HA ha723(p4111,p4115,p4144,p4145);
FA fa1349(p4119,p4123,p3958,p4146,p4147);
HA ha724(p3960,p3964,p4148,p4149);
FA fa1350(p3984,p3988,p4117,p4150,p4151);
HA ha725(p4121,p4125,p4152,p4153);
HA ha726(p4127,p4129,p4154,p4155);
HA ha727(p4133,p4139,p4156,p4157);
HA ha728(p4143,p4145,p4158,p4159);
HA ha729(p3966,p3970,p4160,p4161);
HA ha730(p3978,p3996,p4162,p4163);
FA fa1351(p4131,p4135,p4137,p4164,p4165);
FA fa1352(p4141,p4147,p4149,p4166,p4167);
HA ha731(p4153,p4155,p4168,p4169);
HA ha732(p4157,p4159,p4170,p4171);
FA fa1353(p3980,p3982,p3986,p4172,p4173);
FA fa1354(p3990,p3992,p3994,p4174,p4175);
FA fa1355(p4008,p4010,p4151,p4176,p4177);
FA fa1356(p4161,p4163,p4169,p4178,p4179);
HA ha733(p4171,p3998,p4180,p4181);
FA fa1357(p4000,p4002,p4165,p4182,p4183);
FA fa1358(p4167,p4004,p4006,p4184,p4185);
HA ha734(p4012,p4014,p4186,p4187);
FA fa1359(p4173,p4175,p4177,p4188,p4189);
FA fa1360(p4179,p4181,p4016,p4190,p4191);
FA fa1361(p4018,p4020,p4022,p4192,p4193);
FA fa1362(p4032,p4183,p4187,p4194,p4195);
FA fa1363(p4024,p4026,p4028,p4196,p4197);
FA fa1364(p4185,p4189,p4191,p4198,p4199);
FA fa1365(p4030,p4034,p4042,p4200,p4201);
HA ha735(p4193,p4195,p4202,p4203);
FA fa1366(p4036,p4044,p4197,p4204,p4205);
FA fa1367(p4199,p4203,p4038,p4206,p4207);
FA fa1368(p4040,p4048,p4201,p4208,p4209);
FA fa1369(p4046,p4205,p4207,p4210,p4211);
FA fa1370(p4050,p4054,p4209,p4212,p4213);
FA fa1371(p4052,p4211,p4213,p4214,p4215);
FA fa1372(p4056,p4215,p4058,p4216,p4217);
HA ha736(p4060,p4217,p4218,p4219);
HA ha737(p4219,p4062,p4220,p4221);
HA ha738(ip_0_55,ip_1_54,p4222,p4223);
FA fa1373(ip_2_53,ip_3_52,ip_4_51,p4224,p4225);
HA ha739(ip_5_50,ip_6_49,p4226,p4227);
FA fa1374(ip_7_48,ip_8_47,ip_9_46,p4228,p4229);
HA ha740(ip_10_45,ip_11_44,p4230,p4231);
HA ha741(ip_12_43,ip_13_42,p4232,p4233);
HA ha742(ip_14_41,ip_15_40,p4234,p4235);
FA fa1375(ip_16_39,ip_17_38,ip_18_37,p4236,p4237);
FA fa1376(ip_19_36,ip_20_35,ip_21_34,p4238,p4239);
FA fa1377(ip_22_33,ip_23_32,ip_24_31,p4240,p4241);
FA fa1378(ip_25_30,ip_26_29,ip_27_28,p4242,p4243);
HA ha743(ip_28_27,ip_29_26,p4244,p4245);
FA fa1379(ip_30_25,ip_31_24,ip_32_23,p4246,p4247);
FA fa1380(ip_33_22,ip_34_21,ip_35_20,p4248,p4249);
FA fa1381(ip_36_19,ip_37_18,ip_38_17,p4250,p4251);
FA fa1382(ip_39_16,ip_40_15,ip_41_14,p4252,p4253);
FA fa1383(ip_42_13,ip_43_12,ip_44_11,p4254,p4255);
HA ha744(ip_45_10,ip_46_9,p4256,p4257);
FA fa1384(ip_47_8,ip_48_7,ip_49_6,p4258,p4259);
FA fa1385(ip_50_5,ip_51_4,ip_52_3,p4260,p4261);
FA fa1386(ip_53_2,ip_54_1,ip_55_0,p4262,p4263);
FA fa1387(p4066,p4068,p4074,p4264,p4265);
FA fa1388(p4078,p4080,p4094,p4266,p4267);
HA ha745(p4098,p4223,p4268,p4269);
FA fa1389(p4227,p4231,p4233,p4270,p4271);
FA fa1390(p4235,p4245,p4257,p4272,p4273);
FA fa1391(p4108,p4112,p4225,p4274,p4275);
FA fa1392(p4229,p4237,p4239,p4276,p4277);
HA ha746(p4241,p4243,p4278,p4279);
FA fa1393(p4247,p4249,p4251,p4280,p4281);
FA fa1394(p4253,p4255,p4259,p4282,p4283);
FA fa1395(p4261,p4263,p4269,p4284,p4285);
HA ha747(p4070,p4072,p4286,p4287);
FA fa1396(p4076,p4082,p4084,p4288,p4289);
HA ha748(p4086,p4088,p4290,p4291);
FA fa1397(p4090,p4092,p4096,p4292,p4293);
FA fa1398(p4100,p4102,p4104,p4294,p4295);
HA ha749(p4106,p4118,p4296,p4297);
FA fa1399(p4122,p4265,p4267,p4298,p4299);
FA fa1400(p4271,p4273,p4279,p4300,p4301);
HA ha750(p4110,p4114,p4302,p4303);
HA ha751(p4128,p4132,p4304,p4305);
FA fa1401(p4138,p4142,p4144,p4306,p4307);
FA fa1402(p4275,p4277,p4281,p4308,p4309);
FA fa1403(p4283,p4285,p4287,p4310,p4311);
HA ha752(p4291,p4297,p4312,p4313);
HA ha753(p4116,p4120,p4314,p4315);
HA ha754(p4124,p4126,p4316,p4317);
HA ha755(p4148,p4152,p4318,p4319);
HA ha756(p4154,p4156,p4320,p4321);
FA fa1404(p4158,p4289,p4293,p4322,p4323);
FA fa1405(p4295,p4299,p4301,p4324,p4325);
FA fa1406(p4303,p4305,p4313,p4326,p4327);
FA fa1407(p4130,p4134,p4136,p4328,p4329);
HA ha757(p4140,p4146,p4330,p4331);
FA fa1408(p4160,p4162,p4168,p4332,p4333);
HA ha758(p4170,p4307,p4334,p4335);
FA fa1409(p4309,p4311,p4315,p4336,p4337);
FA fa1410(p4317,p4319,p4321,p4338,p4339);
HA ha759(p4150,p4323,p4340,p4341);
FA fa1411(p4325,p4327,p4331,p4342,p4343);
FA fa1412(p4335,p4164,p4166,p4344,p4345);
FA fa1413(p4180,p4329,p4333,p4346,p4347);
FA fa1414(p4337,p4339,p4341,p4348,p4349);
HA ha760(p4172,p4174,p4350,p4351);
HA ha761(p4176,p4178,p4352,p4353);
FA fa1415(p4186,p4343,p4182,p4354,p4355);
FA fa1416(p4345,p4347,p4349,p4356,p4357);
FA fa1417(p4351,p4353,p4184,p4358,p4359);
HA ha762(p4188,p4190,p4360,p4361);
HA ha763(p4355,p4192,p4362,p4363);
FA fa1418(p4194,p4202,p4357,p4364,p4365);
HA ha764(p4359,p4361,p4366,p4367);
FA fa1419(p4196,p4198,p4363,p4368,p4369);
FA fa1420(p4367,p4200,p4365,p4370,p4371);
FA fa1421(p4204,p4206,p4369,p4372,p4373);
FA fa1422(p4208,p4371,p4210,p4374,p4375);
FA fa1423(p4373,p4212,p4375,p4376,p4377);
FA fa1424(p4214,p4377,p4216,p4378,p4379);
FA fa1425(p4218,p4379,p4220,p4380,p4381);
HA ha765(ip_0_56,ip_1_55,p4382,p4383);
FA fa1426(ip_2_54,ip_3_53,ip_4_52,p4384,p4385);
HA ha766(ip_5_51,ip_6_50,p4386,p4387);
FA fa1427(ip_7_49,ip_8_48,ip_9_47,p4388,p4389);
HA ha767(ip_10_46,ip_11_45,p4390,p4391);
FA fa1428(ip_12_44,ip_13_43,ip_14_42,p4392,p4393);
FA fa1429(ip_15_41,ip_16_40,ip_17_39,p4394,p4395);
HA ha768(ip_18_38,ip_19_37,p4396,p4397);
FA fa1430(ip_20_36,ip_21_35,ip_22_34,p4398,p4399);
FA fa1431(ip_23_33,ip_24_32,ip_25_31,p4400,p4401);
HA ha769(ip_26_30,ip_27_29,p4402,p4403);
FA fa1432(ip_28_28,ip_29_27,ip_30_26,p4404,p4405);
FA fa1433(ip_31_25,ip_32_24,ip_33_23,p4406,p4407);
FA fa1434(ip_34_22,ip_35_21,ip_36_20,p4408,p4409);
HA ha770(ip_37_19,ip_38_18,p4410,p4411);
HA ha771(ip_39_17,ip_40_16,p4412,p4413);
HA ha772(ip_41_15,ip_42_14,p4414,p4415);
FA fa1435(ip_43_13,ip_44_12,ip_45_11,p4416,p4417);
FA fa1436(ip_46_10,ip_47_9,ip_48_8,p4418,p4419);
FA fa1437(ip_49_7,ip_50_6,ip_51_5,p4420,p4421);
HA ha773(ip_52_4,ip_53_3,p4422,p4423);
FA fa1438(ip_54_2,ip_55_1,ip_56_0,p4424,p4425);
HA ha774(p4222,p4226,p4426,p4427);
FA fa1439(p4230,p4232,p4234,p4428,p4429);
HA ha775(p4244,p4256,p4430,p4431);
HA ha776(p4383,p4387,p4432,p4433);
FA fa1440(p4391,p4397,p4403,p4434,p4435);
HA ha777(p4411,p4413,p4436,p4437);
FA fa1441(p4415,p4423,p4268,p4438,p4439);
FA fa1442(p4385,p4389,p4393,p4440,p4441);
FA fa1443(p4395,p4399,p4401,p4442,p4443);
FA fa1444(p4405,p4407,p4409,p4444,p4445);
FA fa1445(p4417,p4419,p4421,p4446,p4447);
FA fa1446(p4425,p4427,p4431,p4448,p4449);
FA fa1447(p4433,p4437,p4224,p4450,p4451);
HA ha778(p4228,p4236,p4452,p4453);
HA ha779(p4238,p4240,p4454,p4455);
HA ha780(p4242,p4246,p4456,p4457);
FA fa1448(p4248,p4250,p4252,p4458,p4459);
FA fa1449(p4254,p4258,p4260,p4460,p4461);
FA fa1450(p4262,p4278,p4429,p4462,p4463);
HA ha781(p4435,p4439,p4464,p4465);
FA fa1451(p4264,p4266,p4270,p4466,p4467);
FA fa1452(p4272,p4286,p4290,p4468,p4469);
FA fa1453(p4296,p4441,p4443,p4470,p4471);
FA fa1454(p4445,p4447,p4449,p4472,p4473);
FA fa1455(p4451,p4453,p4455,p4474,p4475);
FA fa1456(p4457,p4465,p4274,p4476,p4477);
FA fa1457(p4276,p4280,p4282,p4478,p4479);
FA fa1458(p4284,p4302,p4304,p4480,p4481);
FA fa1459(p4312,p4459,p4461,p4482,p4483);
HA ha782(p4463,p4288,p4484,p4485);
HA ha783(p4292,p4294,p4486,p4487);
HA ha784(p4298,p4300,p4488,p4489);
FA fa1460(p4314,p4316,p4318,p4490,p4491);
FA fa1461(p4320,p4467,p4469,p4492,p4493);
FA fa1462(p4471,p4473,p4475,p4494,p4495);
FA fa1463(p4477,p4306,p4308,p4496,p4497);
HA ha785(p4310,p4330,p4498,p4499);
FA fa1464(p4334,p4479,p4481,p4500,p4501);
FA fa1465(p4483,p4485,p4487,p4502,p4503);
FA fa1466(p4489,p4322,p4324,p4504,p4505);
HA ha786(p4326,p4340,p4506,p4507);
FA fa1467(p4491,p4493,p4495,p4508,p4509);
HA ha787(p4499,p4328,p4510,p4511);
FA fa1468(p4332,p4336,p4338,p4512,p4513);
HA ha788(p4497,p4501,p4514,p4515);
FA fa1469(p4503,p4507,p4342,p4516,p4517);
FA fa1470(p4350,p4352,p4505,p4518,p4519);
FA fa1471(p4509,p4511,p4515,p4520,p4521);
FA fa1472(p4344,p4346,p4348,p4522,p4523);
HA ha789(p4513,p4517,p4524,p4525);
HA ha790(p4354,p4360,p4526,p4527);
FA fa1473(p4519,p4521,p4525,p4528,p4529);
HA ha791(p4356,p4358,p4530,p4531);
HA ha792(p4362,p4366,p4532,p4533);
FA fa1474(p4523,p4527,p4529,p4534,p4535);
FA fa1475(p4531,p4533,p4364,p4536,p4537);
FA fa1476(p4535,p4368,p4537,p4538,p4539);
FA fa1477(p4370,p4372,p4539,p4540,p4541);
HA ha793(p4374,p4541,p4542,p4543);
HA ha794(p4376,p4543,p4544,p4545);
HA ha795(p4545,p4378,p4546,p4547);
HA ha796(ip_0_57,ip_1_56,p4548,p4549);
FA fa1478(ip_2_55,ip_3_54,ip_4_53,p4550,p4551);
HA ha797(ip_5_52,ip_6_51,p4552,p4553);
FA fa1479(ip_7_50,ip_8_49,ip_9_48,p4554,p4555);
FA fa1480(ip_10_47,ip_11_46,ip_12_45,p4556,p4557);
HA ha798(ip_13_44,ip_14_43,p4558,p4559);
HA ha799(ip_15_42,ip_16_41,p4560,p4561);
FA fa1481(ip_17_40,ip_18_39,ip_19_38,p4562,p4563);
FA fa1482(ip_20_37,ip_21_36,ip_22_35,p4564,p4565);
FA fa1483(ip_23_34,ip_24_33,ip_25_32,p4566,p4567);
FA fa1484(ip_26_31,ip_27_30,ip_28_29,p4568,p4569);
HA ha800(ip_29_28,ip_30_27,p4570,p4571);
FA fa1485(ip_31_26,ip_32_25,ip_33_24,p4572,p4573);
FA fa1486(ip_34_23,ip_35_22,ip_36_21,p4574,p4575);
FA fa1487(ip_37_20,ip_38_19,ip_39_18,p4576,p4577);
FA fa1488(ip_40_17,ip_41_16,ip_42_15,p4578,p4579);
FA fa1489(ip_43_14,ip_44_13,ip_45_12,p4580,p4581);
HA ha801(ip_46_11,ip_47_10,p4582,p4583);
FA fa1490(ip_48_9,ip_49_8,ip_50_7,p4584,p4585);
FA fa1491(ip_51_6,ip_52_5,ip_53_4,p4586,p4587);
FA fa1492(ip_54_3,ip_55_2,ip_56_1,p4588,p4589);
FA fa1493(ip_57_0,p4382,p4386,p4590,p4591);
FA fa1494(p4390,p4396,p4402,p4592,p4593);
HA ha802(p4410,p4412,p4594,p4595);
HA ha803(p4414,p4422,p4596,p4597);
HA ha804(p4549,p4553,p4598,p4599);
FA fa1495(p4559,p4561,p4571,p4600,p4601);
HA ha805(p4583,p4426,p4602,p4603);
HA ha806(p4430,p4432,p4604,p4605);
FA fa1496(p4436,p4551,p4555,p4606,p4607);
FA fa1497(p4557,p4563,p4565,p4608,p4609);
FA fa1498(p4567,p4569,p4573,p4610,p4611);
HA ha807(p4575,p4577,p4612,p4613);
FA fa1499(p4579,p4581,p4585,p4614,p4615);
FA fa1500(p4587,p4589,p4595,p4616,p4617);
HA ha808(p4597,p4599,p4618,p4619);
HA ha809(p4384,p4388,p4620,p4621);
HA ha810(p4392,p4394,p4622,p4623);
HA ha811(p4398,p4400,p4624,p4625);
HA ha812(p4404,p4406,p4626,p4627);
FA fa1501(p4408,p4416,p4418,p4628,p4629);
HA ha813(p4420,p4424,p4630,p4631);
HA ha814(p4591,p4593,p4632,p4633);
FA fa1502(p4601,p4603,p4605,p4634,p4635);
FA fa1503(p4613,p4619,p4428,p4636,p4637);
HA ha815(p4434,p4438,p4638,p4639);
HA ha816(p4452,p4454,p4640,p4641);
FA fa1504(p4456,p4464,p4607,p4642,p4643);
FA fa1505(p4609,p4611,p4615,p4644,p4645);
HA ha817(p4617,p4621,p4646,p4647);
FA fa1506(p4623,p4625,p4627,p4648,p4649);
HA ha818(p4631,p4633,p4650,p4651);
FA fa1507(p4440,p4442,p4444,p4652,p4653);
HA ha819(p4446,p4448,p4654,p4655);
FA fa1508(p4450,p4629,p4635,p4656,p4657);
FA fa1509(p4637,p4639,p4641,p4658,p4659);
FA fa1510(p4647,p4651,p4458,p4660,p4661);
FA fa1511(p4460,p4462,p4643,p4662,p4663);
FA fa1512(p4645,p4649,p4655,p4664,p4665);
HA ha820(p4466,p4468,p4666,p4667);
HA ha821(p4470,p4472,p4668,p4669);
FA fa1513(p4474,p4476,p4484,p4670,p4671);
FA fa1514(p4486,p4488,p4653,p4672,p4673);
HA ha822(p4657,p4659,p4674,p4675);
FA fa1515(p4661,p4478,p4480,p4676,p4677);
FA fa1516(p4482,p4498,p4663,p4678,p4679);
FA fa1517(p4665,p4667,p4669,p4680,p4681);
FA fa1518(p4675,p4490,p4492,p4682,p4683);
FA fa1519(p4494,p4506,p4671,p4684,p4685);
HA ha823(p4673,p4496,p4686,p4687);
HA ha824(p4500,p4502,p4688,p4689);
HA ha825(p4510,p4514,p4690,p4691);
HA ha826(p4677,p4679,p4692,p4693);
HA ha827(p4681,p4504,p4694,p4695);
HA ha828(p4508,p4683,p4696,p4697);
HA ha829(p4685,p4687,p4698,p4699);
FA fa1520(p4689,p4691,p4693,p4700,p4701);
FA fa1521(p4512,p4516,p4524,p4702,p4703);
FA fa1522(p4695,p4697,p4699,p4704,p4705);
FA fa1523(p4518,p4520,p4526,p4706,p4707);
FA fa1524(p4701,p4522,p4530,p4708,p4709);
FA fa1525(p4532,p4703,p4705,p4710,p4711);
FA fa1526(p4528,p4707,p4534,p4712,p4713);
FA fa1527(p4709,p4711,p4536,p4714,p4715);
HA ha830(p4713,p4715,p4716,p4717);
FA fa1528(p4538,p4717,p4540,p4718,p4719);
FA fa1529(p4542,p4544,p4719,p4720,p4721);
FA fa1530(ip_0_58,ip_1_57,ip_2_56,p4722,p4723);
FA fa1531(ip_3_55,ip_4_54,ip_5_53,p4724,p4725);
FA fa1532(ip_6_52,ip_7_51,ip_8_50,p4726,p4727);
FA fa1533(ip_9_49,ip_10_48,ip_11_47,p4728,p4729);
HA ha831(ip_12_46,ip_13_45,p4730,p4731);
HA ha832(ip_14_44,ip_15_43,p4732,p4733);
HA ha833(ip_16_42,ip_17_41,p4734,p4735);
FA fa1534(ip_18_40,ip_19_39,ip_20_38,p4736,p4737);
FA fa1535(ip_21_37,ip_22_36,ip_23_35,p4738,p4739);
HA ha834(ip_24_34,ip_25_33,p4740,p4741);
FA fa1536(ip_26_32,ip_27_31,ip_28_30,p4742,p4743);
HA ha835(ip_29_29,ip_30_28,p4744,p4745);
FA fa1537(ip_31_27,ip_32_26,ip_33_25,p4746,p4747);
FA fa1538(ip_34_24,ip_35_23,ip_36_22,p4748,p4749);
HA ha836(ip_37_21,ip_38_20,p4750,p4751);
FA fa1539(ip_39_19,ip_40_18,ip_41_17,p4752,p4753);
FA fa1540(ip_42_16,ip_43_15,ip_44_14,p4754,p4755);
FA fa1541(ip_45_13,ip_46_12,ip_47_11,p4756,p4757);
FA fa1542(ip_48_10,ip_49_9,ip_50_8,p4758,p4759);
FA fa1543(ip_51_7,ip_52_6,ip_53_5,p4760,p4761);
HA ha837(ip_54_4,ip_55_3,p4762,p4763);
FA fa1544(ip_56_2,ip_57_1,ip_58_0,p4764,p4765);
FA fa1545(p4548,p4552,p4558,p4766,p4767);
FA fa1546(p4560,p4570,p4582,p4768,p4769);
HA ha838(p4731,p4733,p4770,p4771);
FA fa1547(p4735,p4741,p4745,p4772,p4773);
FA fa1548(p4751,p4763,p4594,p4774,p4775);
HA ha839(p4596,p4598,p4776,p4777);
HA ha840(p4723,p4725,p4778,p4779);
FA fa1549(p4727,p4729,p4737,p4780,p4781);
HA ha841(p4739,p4743,p4782,p4783);
HA ha842(p4747,p4749,p4784,p4785);
FA fa1550(p4753,p4755,p4757,p4786,p4787);
FA fa1551(p4759,p4761,p4765,p4788,p4789);
FA fa1552(p4771,p4550,p4554,p4790,p4791);
FA fa1553(p4556,p4562,p4564,p4792,p4793);
HA ha843(p4566,p4568,p4794,p4795);
HA ha844(p4572,p4574,p4796,p4797);
FA fa1554(p4576,p4578,p4580,p4798,p4799);
FA fa1555(p4584,p4586,p4588,p4800,p4801);
HA ha845(p4602,p4604,p4802,p4803);
HA ha846(p4612,p4618,p4804,p4805);
HA ha847(p4767,p4769,p4806,p4807);
HA ha848(p4773,p4775,p4808,p4809);
FA fa1556(p4777,p4779,p4783,p4810,p4811);
FA fa1557(p4785,p4590,p4592,p4812,p4813);
FA fa1558(p4600,p4620,p4622,p4814,p4815);
HA ha849(p4624,p4626,p4816,p4817);
HA ha850(p4630,p4632,p4818,p4819);
HA ha851(p4781,p4787,p4820,p4821);
HA ha852(p4789,p4795,p4822,p4823);
HA ha853(p4797,p4803,p4824,p4825);
FA fa1559(p4805,p4807,p4809,p4826,p4827);
HA ha854(p4606,p4608,p4828,p4829);
FA fa1560(p4610,p4614,p4616,p4830,p4831);
HA ha855(p4638,p4640,p4832,p4833);
FA fa1561(p4646,p4650,p4791,p4834,p4835);
FA fa1562(p4793,p4799,p4801,p4836,p4837);
FA fa1563(p4811,p4817,p4819,p4838,p4839);
FA fa1564(p4821,p4823,p4825,p4840,p4841);
FA fa1565(p4628,p4634,p4636,p4842,p4843);
FA fa1566(p4654,p4813,p4815,p4844,p4845);
HA ha856(p4827,p4829,p4846,p4847);
FA fa1567(p4833,p4642,p4644,p4848,p4849);
FA fa1568(p4648,p4831,p4835,p4850,p4851);
FA fa1569(p4837,p4839,p4841,p4852,p4853);
FA fa1570(p4847,p4652,p4656,p4854,p4855);
FA fa1571(p4658,p4660,p4666,p4856,p4857);
HA ha857(p4668,p4674,p4858,p4859);
HA ha858(p4843,p4845,p4860,p4861);
HA ha859(p4662,p4664,p4862,p4863);
FA fa1572(p4849,p4851,p4853,p4864,p4865);
HA ha860(p4859,p4861,p4866,p4867);
FA fa1573(p4670,p4672,p4855,p4868,p4869);
HA ha861(p4857,p4863,p4870,p4871);
FA fa1574(p4867,p4676,p4678,p4872,p4873);
FA fa1575(p4680,p4686,p4688,p4874,p4875);
HA ha862(p4690,p4692,p4876,p4877);
HA ha863(p4865,p4871,p4878,p4879);
FA fa1576(p4682,p4684,p4694,p4880,p4881);
FA fa1577(p4696,p4698,p4869,p4882,p4883);
FA fa1578(p4877,p4879,p4873,p4884,p4885);
HA ha864(p4875,p4700,p4886,p4887);
FA fa1579(p4881,p4883,p4885,p4888,p4889);
HA ha865(p4702,p4704,p4890,p4891);
FA fa1580(p4887,p4706,p4889,p4892,p4893);
FA fa1581(p4891,p4708,p4710,p4894,p4895);
FA fa1582(p4712,p4893,p4714,p4896,p4897);
FA fa1583(p4716,p4895,p4897,p4898,p4899);
HA ha866(p4899,p4718,p4900,p4901);
FA fa1584(ip_0_59,ip_1_58,ip_2_57,p4902,p4903);
FA fa1585(ip_3_56,ip_4_55,ip_5_54,p4904,p4905);
FA fa1586(ip_6_53,ip_7_52,ip_8_51,p4906,p4907);
HA ha867(ip_9_50,ip_10_49,p4908,p4909);
FA fa1587(ip_11_48,ip_12_47,ip_13_46,p4910,p4911);
HA ha868(ip_14_45,ip_15_44,p4912,p4913);
HA ha869(ip_16_43,ip_17_42,p4914,p4915);
HA ha870(ip_18_41,ip_19_40,p4916,p4917);
FA fa1588(ip_20_39,ip_21_38,ip_22_37,p4918,p4919);
FA fa1589(ip_23_36,ip_24_35,ip_25_34,p4920,p4921);
FA fa1590(ip_26_33,ip_27_32,ip_28_31,p4922,p4923);
HA ha871(ip_29_30,ip_30_29,p4924,p4925);
FA fa1591(ip_31_28,ip_32_27,ip_33_26,p4926,p4927);
HA ha872(ip_34_25,ip_35_24,p4928,p4929);
FA fa1592(ip_36_23,ip_37_22,ip_38_21,p4930,p4931);
FA fa1593(ip_39_20,ip_40_19,ip_41_18,p4932,p4933);
FA fa1594(ip_42_17,ip_43_16,ip_44_15,p4934,p4935);
FA fa1595(ip_45_14,ip_46_13,ip_47_12,p4936,p4937);
FA fa1596(ip_48_11,ip_49_10,ip_50_9,p4938,p4939);
FA fa1597(ip_51_8,ip_52_7,ip_53_6,p4940,p4941);
FA fa1598(ip_54_5,ip_55_4,ip_56_3,p4942,p4943);
HA ha873(ip_57_2,ip_58_1,p4944,p4945);
HA ha874(ip_59_0,p4730,p4946,p4947);
HA ha875(p4732,p4734,p4948,p4949);
FA fa1599(p4740,p4744,p4750,p4950,p4951);
FA fa1600(p4762,p4909,p4913,p4952,p4953);
FA fa1601(p4915,p4917,p4925,p4954,p4955);
FA fa1602(p4929,p4945,p4770,p4956,p4957);
HA ha876(p4903,p4905,p4958,p4959);
HA ha877(p4907,p4911,p4960,p4961);
FA fa1603(p4919,p4921,p4923,p4962,p4963);
FA fa1604(p4927,p4931,p4933,p4964,p4965);
FA fa1605(p4935,p4937,p4939,p4966,p4967);
FA fa1606(p4941,p4943,p4947,p4968,p4969);
FA fa1607(p4949,p4722,p4724,p4970,p4971);
FA fa1608(p4726,p4728,p4736,p4972,p4973);
FA fa1609(p4738,p4742,p4746,p4974,p4975);
HA ha878(p4748,p4752,p4976,p4977);
HA ha879(p4754,p4756,p4978,p4979);
HA ha880(p4758,p4760,p4980,p4981);
HA ha881(p4764,p4776,p4982,p4983);
HA ha882(p4778,p4782,p4984,p4985);
HA ha883(p4784,p4951,p4986,p4987);
FA fa1610(p4953,p4955,p4957,p4988,p4989);
FA fa1611(p4959,p4961,p4766,p4990,p4991);
HA ha884(p4768,p4772,p4992,p4993);
FA fa1612(p4774,p4794,p4796,p4994,p4995);
HA ha885(p4802,p4804,p4996,p4997);
FA fa1613(p4806,p4808,p4963,p4998,p4999);
FA fa1614(p4965,p4967,p4969,p5000,p5001);
HA ha886(p4977,p4979,p5002,p5003);
FA fa1615(p4981,p4983,p4985,p5004,p5005);
FA fa1616(p4987,p4780,p4786,p5006,p5007);
HA ha887(p4788,p4816,p5008,p5009);
HA ha888(p4818,p4820,p5010,p5011);
FA fa1617(p4822,p4824,p4971,p5012,p5013);
HA ha889(p4973,p4975,p5014,p5015);
FA fa1618(p4989,p4991,p4993,p5016,p5017);
FA fa1619(p4997,p5003,p4790,p5018,p5019);
FA fa1620(p4792,p4798,p4800,p5020,p5021);
HA ha890(p4810,p4828,p5022,p5023);
HA ha891(p4832,p4995,p5024,p5025);
FA fa1621(p4999,p5001,p5005,p5026,p5027);
HA ha892(p5009,p5011,p5028,p5029);
FA fa1622(p5015,p4812,p4814,p5030,p5031);
HA ha893(p4826,p4846,p5032,p5033);
FA fa1623(p5007,p5013,p5017,p5034,p5035);
HA ha894(p5019,p5023,p5036,p5037);
HA ha895(p5025,p5029,p5038,p5039);
HA ha896(p4830,p4834,p5040,p5041);
HA ha897(p4836,p4838,p5042,p5043);
HA ha898(p4840,p5021,p5044,p5045);
FA fa1624(p5027,p5033,p5037,p5046,p5047);
FA fa1625(p5039,p4842,p4844,p5048,p5049);
HA ha899(p4858,p4860,p5050,p5051);
HA ha900(p5031,p5035,p5052,p5053);
FA fa1626(p5041,p5043,p5045,p5054,p5055);
HA ha901(p4848,p4850,p5056,p5057);
FA fa1627(p4852,p4862,p4866,p5058,p5059);
HA ha902(p5047,p5051,p5060,p5061);
FA fa1628(p5053,p4854,p4856,p5062,p5063);
HA ha903(p4870,p5049,p5064,p5065);
HA ha904(p5055,p5057,p5066,p5067);
FA fa1629(p5061,p4864,p4876,p5068,p5069);
FA fa1630(p4878,p5059,p5065,p5070,p5071);
FA fa1631(p5067,p4868,p5063,p5072,p5073);
FA fa1632(p4872,p4874,p5069,p5074,p5075);
FA fa1633(p5071,p4880,p4882,p5076,p5077);
FA fa1634(p4884,p4886,p5073,p5078,p5079);
FA fa1635(p4890,p5075,p4888,p5080,p5081);
FA fa1636(p5077,p5079,p5081,p5082,p5083);
HA ha905(p4892,p5083,p5084,p5085);
FA fa1637(p4894,p5085,p4896,p5086,p5087);
FA fa1638(p4898,p5087,p4900,p5088,p5089);
HA ha906(ip_0_60,ip_1_59,p5090,p5091);
FA fa1639(ip_2_58,ip_3_57,ip_4_56,p5092,p5093);
FA fa1640(ip_5_55,ip_6_54,ip_7_53,p5094,p5095);
FA fa1641(ip_8_52,ip_9_51,ip_10_50,p5096,p5097);
HA ha907(ip_11_49,ip_12_48,p5098,p5099);
HA ha908(ip_13_47,ip_14_46,p5100,p5101);
FA fa1642(ip_15_45,ip_16_44,ip_17_43,p5102,p5103);
HA ha909(ip_18_42,ip_19_41,p5104,p5105);
FA fa1643(ip_20_40,ip_21_39,ip_22_38,p5106,p5107);
FA fa1644(ip_23_37,ip_24_36,ip_25_35,p5108,p5109);
HA ha910(ip_26_34,ip_27_33,p5110,p5111);
FA fa1645(ip_28_32,ip_29_31,ip_30_30,p5112,p5113);
FA fa1646(ip_31_29,ip_32_28,ip_33_27,p5114,p5115);
FA fa1647(ip_34_26,ip_35_25,ip_36_24,p5116,p5117);
FA fa1648(ip_37_23,ip_38_22,ip_39_21,p5118,p5119);
HA ha911(ip_40_20,ip_41_19,p5120,p5121);
FA fa1649(ip_42_18,ip_43_17,ip_44_16,p5122,p5123);
FA fa1650(ip_45_15,ip_46_14,ip_47_13,p5124,p5125);
HA ha912(ip_48_12,ip_49_11,p5126,p5127);
HA ha913(ip_50_10,ip_51_9,p5128,p5129);
FA fa1651(ip_52_8,ip_53_7,ip_54_6,p5130,p5131);
FA fa1652(ip_55_5,ip_56_4,ip_57_3,p5132,p5133);
FA fa1653(ip_58_2,ip_59_1,ip_60_0,p5134,p5135);
FA fa1654(p4908,p4912,p4914,p5136,p5137);
FA fa1655(p4916,p4924,p4928,p5138,p5139);
HA ha914(p4944,p5091,p5140,p5141);
HA ha915(p5099,p5101,p5142,p5143);
HA ha916(p5105,p5111,p5144,p5145);
HA ha917(p5121,p5127,p5146,p5147);
HA ha918(p5129,p4946,p5148,p5149);
FA fa1656(p4948,p5093,p5095,p5150,p5151);
HA ha919(p5097,p5103,p5152,p5153);
FA fa1657(p5107,p5109,p5113,p5154,p5155);
HA ha920(p5115,p5117,p5156,p5157);
FA fa1658(p5119,p5123,p5125,p5158,p5159);
FA fa1659(p5131,p5133,p5135,p5160,p5161);
FA fa1660(p5141,p5143,p5145,p5162,p5163);
HA ha921(p5147,p4902,p5164,p5165);
HA ha922(p4904,p4906,p5166,p5167);
FA fa1661(p4910,p4918,p4920,p5168,p5169);
FA fa1662(p4922,p4926,p4930,p5170,p5171);
HA ha923(p4932,p4934,p5172,p5173);
HA ha924(p4936,p4938,p5174,p5175);
HA ha925(p4940,p4942,p5176,p5177);
FA fa1663(p4958,p4960,p5137,p5178,p5179);
FA fa1664(p5139,p5149,p5153,p5180,p5181);
FA fa1665(p5157,p4950,p4952,p5182,p5183);
FA fa1666(p4954,p4956,p4976,p5184,p5185);
HA ha926(p4978,p4980,p5186,p5187);
HA ha927(p4982,p4984,p5188,p5189);
FA fa1667(p4986,p5151,p5155,p5190,p5191);
FA fa1668(p5159,p5161,p5163,p5192,p5193);
HA ha928(p5165,p5167,p5194,p5195);
FA fa1669(p5173,p5175,p5177,p5196,p5197);
HA ha929(p4962,p4964,p5198,p5199);
FA fa1670(p4966,p4968,p4992,p5200,p5201);
FA fa1671(p4996,p5002,p5169,p5202,p5203);
HA ha930(p5171,p5179,p5204,p5205);
HA ha931(p5181,p5187,p5206,p5207);
HA ha932(p5189,p5195,p5208,p5209);
FA fa1672(p4970,p4972,p4974,p5210,p5211);
HA ha933(p4988,p4990,p5212,p5213);
FA fa1673(p5008,p5010,p5014,p5214,p5215);
HA ha934(p5183,p5185,p5216,p5217);
FA fa1674(p5191,p5193,p5197,p5218,p5219);
HA ha935(p5199,p5205,p5220,p5221);
FA fa1675(p5207,p5209,p4994,p5222,p5223);
FA fa1676(p4998,p5000,p5004,p5224,p5225);
FA fa1677(p5022,p5024,p5028,p5226,p5227);
HA ha936(p5201,p5203,p5228,p5229);
HA ha937(p5213,p5217,p5230,p5231);
FA fa1678(p5221,p5006,p5012,p5232,p5233);
HA ha938(p5016,p5018,p5234,p5235);
HA ha939(p5032,p5036,p5236,p5237);
HA ha940(p5038,p5211,p5238,p5239);
FA fa1679(p5215,p5219,p5223,p5240,p5241);
HA ha941(p5229,p5231,p5242,p5243);
HA ha942(p5020,p5026,p5244,p5245);
HA ha943(p5040,p5042,p5246,p5247);
HA ha944(p5044,p5225,p5248,p5249);
HA ha945(p5227,p5235,p5250,p5251);
FA fa1680(p5237,p5239,p5243,p5252,p5253);
HA ha946(p5030,p5034,p5254,p5255);
FA fa1681(p5050,p5052,p5233,p5256,p5257);
FA fa1682(p5241,p5245,p5247,p5258,p5259);
FA fa1683(p5249,p5251,p5046,p5260,p5261);
FA fa1684(p5056,p5060,p5253,p5262,p5263);
FA fa1685(p5255,p5048,p5054,p5264,p5265);
FA fa1686(p5064,p5066,p5257,p5266,p5267);
HA ha947(p5259,p5261,p5268,p5269);
HA ha948(p5058,p5263,p5270,p5271);
FA fa1687(p5269,p5062,p5265,p5272,p5273);
HA ha949(p5267,p5271,p5274,p5275);
FA fa1688(p5068,p5070,p5275,p5276,p5277);
FA fa1689(p5072,p5273,p5074,p5278,p5279);
HA ha950(p5277,p5076,p5280,p5281);
FA fa1690(p5078,p5279,p5080,p5282,p5283);
HA ha951(p5281,p5082,p5284,p5285);
FA fa1691(p5084,p5283,p5285,p5286,p5287);
HA ha952(p5287,p5086,p5288,p5289);
FA fa1692(ip_0_61,ip_1_60,ip_2_59,p5290,p5291);
FA fa1693(ip_3_58,ip_4_57,ip_5_56,p5292,p5293);
FA fa1694(ip_6_55,ip_7_54,ip_8_53,p5294,p5295);
HA ha953(ip_9_52,ip_10_51,p5296,p5297);
HA ha954(ip_11_50,ip_12_49,p5298,p5299);
FA fa1695(ip_13_48,ip_14_47,ip_15_46,p5300,p5301);
HA ha955(ip_16_45,ip_17_44,p5302,p5303);
FA fa1696(ip_18_43,ip_19_42,ip_20_41,p5304,p5305);
FA fa1697(ip_21_40,ip_22_39,ip_23_38,p5306,p5307);
FA fa1698(ip_24_37,ip_25_36,ip_26_35,p5308,p5309);
FA fa1699(ip_27_34,ip_28_33,ip_29_32,p5310,p5311);
FA fa1700(ip_30_31,ip_31_30,ip_32_29,p5312,p5313);
FA fa1701(ip_33_28,ip_34_27,ip_35_26,p5314,p5315);
HA ha956(ip_36_25,ip_37_24,p5316,p5317);
FA fa1702(ip_38_23,ip_39_22,ip_40_21,p5318,p5319);
FA fa1703(ip_41_20,ip_42_19,ip_43_18,p5320,p5321);
FA fa1704(ip_44_17,ip_45_16,ip_46_15,p5322,p5323);
FA fa1705(ip_47_14,ip_48_13,ip_49_12,p5324,p5325);
FA fa1706(ip_50_11,ip_51_10,ip_52_9,p5326,p5327);
HA ha957(ip_53_8,ip_54_7,p5328,p5329);
FA fa1707(ip_55_6,ip_56_5,ip_57_4,p5330,p5331);
FA fa1708(ip_58_3,ip_59_2,ip_60_1,p5332,p5333);
FA fa1709(ip_61_0,p5090,p5098,p5334,p5335);
HA ha958(p5100,p5104,p5336,p5337);
FA fa1710(p5110,p5120,p5126,p5338,p5339);
FA fa1711(p5128,p5297,p5299,p5340,p5341);
FA fa1712(p5303,p5317,p5329,p5342,p5343);
FA fa1713(p5140,p5142,p5144,p5344,p5345);
FA fa1714(p5146,p5291,p5293,p5346,p5347);
FA fa1715(p5295,p5301,p5305,p5348,p5349);
FA fa1716(p5307,p5309,p5311,p5350,p5351);
HA ha959(p5313,p5315,p5352,p5353);
HA ha960(p5319,p5321,p5354,p5355);
HA ha961(p5323,p5325,p5356,p5357);
FA fa1717(p5327,p5331,p5333,p5358,p5359);
HA ha962(p5337,p5092,p5360,p5361);
HA ha963(p5094,p5096,p5362,p5363);
HA ha964(p5102,p5106,p5364,p5365);
FA fa1718(p5108,p5112,p5114,p5366,p5367);
HA ha965(p5116,p5118,p5368,p5369);
FA fa1719(p5122,p5124,p5130,p5370,p5371);
FA fa1720(p5132,p5134,p5148,p5372,p5373);
FA fa1721(p5152,p5156,p5335,p5374,p5375);
FA fa1722(p5339,p5341,p5343,p5376,p5377);
FA fa1723(p5353,p5355,p5357,p5378,p5379);
HA ha966(p5136,p5138,p5380,p5381);
FA fa1724(p5164,p5166,p5172,p5382,p5383);
FA fa1725(p5174,p5176,p5345,p5384,p5385);
FA fa1726(p5347,p5349,p5351,p5386,p5387);
HA ha967(p5359,p5361,p5388,p5389);
HA ha968(p5363,p5365,p5390,p5391);
HA ha969(p5369,p5150,p5392,p5393);
HA ha970(p5154,p5158,p5394,p5395);
HA ha971(p5160,p5162,p5396,p5397);
HA ha972(p5186,p5188,p5398,p5399);
FA fa1727(p5194,p5367,p5371,p5400,p5401);
HA ha973(p5373,p5375,p5402,p5403);
HA ha974(p5377,p5379,p5404,p5405);
FA fa1728(p5381,p5389,p5391,p5406,p5407);
HA ha975(p5168,p5170,p5408,p5409);
HA ha976(p5178,p5180,p5410,p5411);
HA ha977(p5198,p5204,p5412,p5413);
FA fa1729(p5206,p5208,p5383,p5414,p5415);
FA fa1730(p5385,p5387,p5393,p5416,p5417);
FA fa1731(p5395,p5397,p5399,p5418,p5419);
HA ha978(p5403,p5405,p5420,p5421);
FA fa1732(p5182,p5184,p5190,p5422,p5423);
FA fa1733(p5192,p5196,p5212,p5424,p5425);
HA ha979(p5216,p5220,p5426,p5427);
FA fa1734(p5401,p5407,p5409,p5428,p5429);
HA ha980(p5411,p5413,p5430,p5431);
FA fa1735(p5421,p5200,p5202,p5432,p5433);
HA ha981(p5228,p5230,p5434,p5435);
FA fa1736(p5415,p5417,p5419,p5436,p5437);
FA fa1737(p5427,p5431,p5210,p5438,p5439);
FA fa1738(p5214,p5218,p5222,p5440,p5441);
HA ha982(p5234,p5236,p5442,p5443);
HA ha983(p5238,p5242,p5444,p5445);
FA fa1739(p5423,p5425,p5429,p5446,p5447);
FA fa1740(p5435,p5224,p5226,p5448,p5449);
HA ha984(p5244,p5246,p5450,p5451);
HA ha985(p5248,p5250,p5452,p5453);
HA ha986(p5433,p5437,p5454,p5455);
FA fa1741(p5439,p5443,p5445,p5456,p5457);
FA fa1742(p5232,p5240,p5254,p5458,p5459);
HA ha987(p5441,p5447,p5460,p5461);
FA fa1743(p5451,p5453,p5455,p5462,p5463);
FA fa1744(p5252,p5449,p5457,p5464,p5465);
FA fa1745(p5461,p5256,p5258,p5466,p5467);
HA ha988(p5260,p5268,p5468,p5469);
FA fa1746(p5459,p5463,p5262,p5470,p5471);
HA ha989(p5270,p5465,p5472,p5473);
HA ha990(p5469,p5264,p5474,p5475);
FA fa1747(p5266,p5274,p5467,p5476,p5477);
FA fa1748(p5471,p5473,p5475,p5478,p5479);
FA fa1749(p5272,p5477,p5479,p5480,p5481);
FA fa1750(p5276,p5278,p5280,p5482,p5483);
FA fa1751(p5481,p5282,p5284,p5484,p5485);
FA fa1752(p5483,p5286,p5485,p5486,p5487);
FA fa1753(ip_0_62,ip_1_61,ip_2_60,p5488,p5489);
FA fa1754(ip_3_59,ip_4_58,ip_5_57,p5490,p5491);
HA ha991(ip_6_56,ip_7_55,p5492,p5493);
HA ha992(ip_8_54,ip_9_53,p5494,p5495);
FA fa1755(ip_10_52,ip_11_51,ip_12_50,p5496,p5497);
FA fa1756(ip_13_49,ip_14_48,ip_15_47,p5498,p5499);
FA fa1757(ip_16_46,ip_17_45,ip_18_44,p5500,p5501);
HA ha993(ip_19_43,ip_20_42,p5502,p5503);
FA fa1758(ip_21_41,ip_22_40,ip_23_39,p5504,p5505);
FA fa1759(ip_24_38,ip_25_37,ip_26_36,p5506,p5507);
HA ha994(ip_27_35,ip_28_34,p5508,p5509);
FA fa1760(ip_29_33,ip_30_32,ip_31_31,p5510,p5511);
HA ha995(ip_32_30,ip_33_29,p5512,p5513);
FA fa1761(ip_34_28,ip_35_27,ip_36_26,p5514,p5515);
FA fa1762(ip_37_25,ip_38_24,ip_39_23,p5516,p5517);
HA ha996(ip_40_22,ip_41_21,p5518,p5519);
HA ha997(ip_42_20,ip_43_19,p5520,p5521);
FA fa1763(ip_44_18,ip_45_17,ip_46_16,p5522,p5523);
HA ha998(ip_47_15,ip_48_14,p5524,p5525);
HA ha999(ip_49_13,ip_50_12,p5526,p5527);
FA fa1764(ip_51_11,ip_52_10,ip_53_9,p5528,p5529);
FA fa1765(ip_54_8,ip_55_7,ip_56_6,p5530,p5531);
HA ha1000(ip_57_5,ip_58_4,p5532,p5533);
FA fa1766(ip_59_3,ip_60_2,ip_61_1,p5534,p5535);
HA ha1001(ip_62_0,p5296,p5536,p5537);
HA ha1002(p5298,p5302,p5538,p5539);
HA ha1003(p5316,p5328,p5540,p5541);
FA fa1767(p5493,p5495,p5503,p5542,p5543);
FA fa1768(p5509,p5513,p5519,p5544,p5545);
FA fa1769(p5521,p5525,p5527,p5546,p5547);
HA ha1004(p5533,p5336,p5548,p5549);
HA ha1005(p5489,p5491,p5550,p5551);
FA fa1770(p5497,p5499,p5501,p5552,p5553);
FA fa1771(p5505,p5507,p5511,p5554,p5555);
FA fa1772(p5515,p5517,p5523,p5556,p5557);
HA ha1006(p5529,p5531,p5558,p5559);
FA fa1773(p5535,p5537,p5539,p5560,p5561);
HA ha1007(p5541,p5290,p5562,p5563);
HA ha1008(p5292,p5294,p5564,p5565);
HA ha1009(p5300,p5304,p5566,p5567);
FA fa1774(p5306,p5308,p5310,p5568,p5569);
FA fa1775(p5312,p5314,p5318,p5570,p5571);
HA ha1010(p5320,p5322,p5572,p5573);
FA fa1776(p5324,p5326,p5330,p5574,p5575);
FA fa1777(p5332,p5352,p5354,p5576,p5577);
FA fa1778(p5356,p5543,p5545,p5578,p5579);
HA ha1011(p5547,p5549,p5580,p5581);
FA fa1779(p5551,p5559,p5334,p5582,p5583);
HA ha1012(p5338,p5340,p5584,p5585);
FA fa1780(p5342,p5360,p5362,p5586,p5587);
FA fa1781(p5364,p5368,p5553,p5588,p5589);
FA fa1782(p5555,p5557,p5561,p5590,p5591);
HA ha1013(p5563,p5565,p5592,p5593);
FA fa1783(p5567,p5573,p5581,p5594,p5595);
FA fa1784(p5344,p5346,p5348,p5596,p5597);
FA fa1785(p5350,p5358,p5380,p5598,p5599);
FA fa1786(p5388,p5390,p5569,p5600,p5601);
FA fa1787(p5571,p5575,p5577,p5602,p5603);
FA fa1788(p5579,p5583,p5585,p5604,p5605);
FA fa1789(p5593,p5366,p5370,p5606,p5607);
FA fa1790(p5372,p5374,p5376,p5608,p5609);
FA fa1791(p5378,p5392,p5394,p5610,p5611);
FA fa1792(p5396,p5398,p5402,p5612,p5613);
FA fa1793(p5404,p5587,p5589,p5614,p5615);
FA fa1794(p5591,p5595,p5382,p5616,p5617);
HA ha1014(p5384,p5386,p5618,p5619);
FA fa1795(p5408,p5410,p5412,p5620,p5621);
HA ha1015(p5420,p5597,p5622,p5623);
HA ha1016(p5599,p5601,p5624,p5625);
FA fa1796(p5603,p5605,p5400,p5626,p5627);
HA ha1017(p5406,p5426,p5628,p5629);
FA fa1797(p5430,p5607,p5609,p5630,p5631);
HA ha1018(p5611,p5613,p5632,p5633);
HA ha1019(p5615,p5617,p5634,p5635);
HA ha1020(p5619,p5623,p5636,p5637);
FA fa1798(p5625,p5414,p5416,p5638,p5639);
HA ha1021(p5418,p5434,p5640,p5641);
HA ha1022(p5621,p5627,p5642,p5643);
FA fa1799(p5629,p5633,p5635,p5644,p5645);
FA fa1800(p5637,p5422,p5424,p5646,p5647);
HA ha1023(p5428,p5442,p5648,p5649);
FA fa1801(p5444,p5631,p5641,p5650,p5651);
HA ha1024(p5643,p5432,p5652,p5653);
FA fa1802(p5436,p5438,p5450,p5654,p5655);
HA ha1025(p5452,p5454,p5656,p5657);
FA fa1803(p5639,p5645,p5649,p5658,p5659);
FA fa1804(p5440,p5446,p5460,p5660,p5661);
HA ha1026(p5647,p5651,p5662,p5663);
FA fa1805(p5653,p5657,p5448,p5664,p5665);
HA ha1027(p5456,p5655,p5666,p5667);
HA ha1028(p5659,p5663,p5668,p5669);
FA fa1806(p5458,p5462,p5468,p5670,p5671);
FA fa1807(p5661,p5665,p5667,p5672,p5673);
HA ha1029(p5669,p5464,p5674,p5675);
FA fa1808(p5472,p5466,p5470,p5676,p5677);
FA fa1809(p5474,p5671,p5673,p5678,p5679);
HA ha1030(p5675,p5476,p5680,p5681);
FA fa1810(p5478,p5677,p5679,p5682,p5683);
HA ha1031(p5681,p5480,p5684,p5685);
FA fa1811(p5683,p5685,p5482,p5686,p5687);
FA fa1812(p5687,p5484,p5486,p5688,p5689);
FA fa1813(ip_0_63,ip_1_62,ip_2_61,p5690,p5691);
FA fa1814(ip_3_60,ip_4_59,ip_5_58,p5692,p5693);
HA ha1032(ip_6_57,ip_7_56,p5694,p5695);
FA fa1815(ip_8_55,ip_9_54,ip_10_53,p5696,p5697);
FA fa1816(ip_11_52,ip_12_51,ip_13_50,p5698,p5699);
FA fa1817(ip_14_49,ip_15_48,ip_16_47,p5700,p5701);
FA fa1818(ip_17_46,ip_18_45,ip_19_44,p5702,p5703);
FA fa1819(ip_20_43,ip_21_42,ip_22_41,p5704,p5705);
FA fa1820(ip_23_40,ip_24_39,ip_25_38,p5706,p5707);
HA ha1033(ip_26_37,ip_27_36,p5708,p5709);
FA fa1821(ip_28_35,ip_29_34,ip_30_33,p5710,p5711);
FA fa1822(ip_31_32,ip_32_31,ip_33_30,p5712,p5713);
HA ha1034(ip_34_29,ip_35_28,p5714,p5715);
FA fa1823(ip_36_27,ip_37_26,ip_38_25,p5716,p5717);
FA fa1824(ip_39_24,ip_40_23,ip_41_22,p5718,p5719);
HA ha1035(ip_42_21,ip_43_20,p5720,p5721);
FA fa1825(ip_44_19,ip_45_18,ip_46_17,p5722,p5723);
FA fa1826(ip_47_16,ip_48_15,ip_49_14,p5724,p5725);
FA fa1827(ip_50_13,ip_51_12,ip_52_11,p5726,p5727);
HA ha1036(ip_53_10,ip_54_9,p5728,p5729);
FA fa1828(ip_55_8,ip_56_7,ip_57_6,p5730,p5731);
HA ha1037(ip_58_5,ip_59_4,p5732,p5733);
HA ha1038(ip_60_3,ip_61_2,p5734,p5735);
FA fa1829(ip_62_1,ip_63_0,p5492,p5736,p5737);
FA fa1830(p5494,p5502,p5508,p5738,p5739);
HA ha1039(p5512,p5518,p5740,p5741);
FA fa1831(p5520,p5524,p5526,p5742,p5743);
FA fa1832(p5532,p5695,p5709,p5744,p5745);
HA ha1040(p5715,p5721,p5746,p5747);
HA ha1041(p5729,p5733,p5748,p5749);
HA ha1042(p5735,p5536,p5750,p5751);
FA fa1833(p5538,p5540,p5691,p5752,p5753);
FA fa1834(p5693,p5697,p5699,p5754,p5755);
HA ha1043(p5701,p5703,p5756,p5757);
FA fa1835(p5705,p5707,p5711,p5758,p5759);
FA fa1836(p5713,p5717,p5719,p5760,p5761);
FA fa1837(p5723,p5725,p5727,p5762,p5763);
HA ha1044(p5731,p5737,p5764,p5765);
FA fa1838(p5741,p5747,p5749,p5766,p5767);
FA fa1839(p5488,p5490,p5496,p5768,p5769);
FA fa1840(p5498,p5500,p5504,p5770,p5771);
FA fa1841(p5506,p5510,p5514,p5772,p5773);
FA fa1842(p5516,p5522,p5528,p5774,p5775);
FA fa1843(p5530,p5534,p5548,p5776,p5777);
FA fa1844(p5550,p5558,p5739,p5778,p5779);
FA fa1845(p5743,p5745,p5751,p5780,p5781);
HA ha1045(p5757,p5765,p5782,p5783);
HA ha1046(p5542,p5544,p5784,p5785);
FA fa1846(p5546,p5562,p5564,p5786,p5787);
HA ha1047(p5566,p5572,p5788,p5789);
HA ha1048(p5580,p5753,p5790,p5791);
FA fa1847(p5755,p5759,p5761,p5792,p5793);
FA fa1848(p5763,p5767,p5783,p5794,p5795);
FA fa1849(p5552,p5554,p5556,p5796,p5797);
HA ha1049(p5560,p5584,p5798,p5799);
FA fa1850(p5592,p5769,p5771,p5800,p5801);
HA ha1050(p5773,p5775,p5802,p5803);
FA fa1851(p5777,p5779,p5781,p5804,p5805);
FA fa1852(p5785,p5789,p5791,p5806,p5807);
FA fa1853(p5568,p5570,p5574,p5808,p5809);
FA fa1854(p5576,p5578,p5582,p5810,p5811);
FA fa1855(p5787,p5793,p5795,p5812,p5813);
FA fa1856(p5799,p5803,p5586,p5814,p5815);
FA fa1857(p5588,p5590,p5594,p5816,p5817);
FA fa1858(p5797,p5801,p5805,p5818,p5819);
FA fa1859(p5807,p5596,p5598,p5820,p5821);
HA ha1051(p5600,p5602,p5822,p5823);
FA fa1860(p5604,p5618,p5622,p5824,p5825);
FA fa1861(p5624,p5809,p5811,p5826,p5827);
HA ha1052(p5813,p5815,p5828,p5829);
FA fa1862(p5606,p5608,p5610,p5830,p5831);
FA fa1863(p5612,p5614,p5616,p5832,p5833);
HA ha1053(p5628,p5632,p5834,p5835);
FA fa1864(p5634,p5636,p5817,p5836,p5837);
HA ha1054(p5819,p5823,p5838,p5839);
HA ha1055(p5829,p5620,p5840,p5841);
FA fa1865(p5626,p5640,p5642,p5842,p5843);
FA fa1866(p5821,p5825,p5827,p5844,p5845);
HA ha1056(p5835,p5839,p5846,p5847);
FA fa1867(p5630,p5648,p5831,p5848,p5849);
FA fa1868(p5833,p5837,p5841,p5850,p5851);
FA fa1869(p5847,p5638,p5644,p5852,p5853);
FA fa1870(p5652,p5656,p5843,p5854,p5855);
FA fa1871(p5845,p5646,p5650,p5856,p5857);
HA ha1057(p5662,p5849,p5858,p5859);
FA fa1872(p5851,p5654,p5658,p5860,p5861);
FA fa1873(p5666,p5668,p5853,p5862,p5863);
HA ha1058(p5855,p5859,p5864,p5865);
FA fa1874(p5660,p5664,p5857,p5866,p5867);
FA fa1875(p5865,p5674,p5861,p5868,p5869);
HA ha1059(p5863,p5670,p5870,p5871);
HA ha1060(p5672,p5867,p5872,p5873);
FA fa1876(p5869,p5871,p5873,p5874,p5875);
FA fa1877(p5676,p5678,p5680,p5876,p5877);
FA fa1878(p5875,p5682,p5684,p5878,p5879);
FA fa1879(p5877,p5879,p5686,p5880,p5881);
FA fa1880(ip_1_63,ip_2_62,ip_3_61,p5882,p5883);
FA fa1881(ip_4_60,ip_5_59,ip_6_58,p5884,p5885);
HA ha1061(ip_7_57,ip_8_56,p5886,p5887);
HA ha1062(ip_9_55,ip_10_54,p5888,p5889);
HA ha1063(ip_11_53,ip_12_52,p5890,p5891);
FA fa1882(ip_13_51,ip_14_50,ip_15_49,p5892,p5893);
FA fa1883(ip_16_48,ip_17_47,ip_18_46,p5894,p5895);
FA fa1884(ip_19_45,ip_20_44,ip_21_43,p5896,p5897);
FA fa1885(ip_22_42,ip_23_41,ip_24_40,p5898,p5899);
HA ha1064(ip_25_39,ip_26_38,p5900,p5901);
FA fa1886(ip_27_37,ip_28_36,ip_29_35,p5902,p5903);
HA ha1065(ip_30_34,ip_31_33,p5904,p5905);
FA fa1887(ip_32_32,ip_33_31,ip_34_30,p5906,p5907);
FA fa1888(ip_35_29,ip_36_28,ip_37_27,p5908,p5909);
FA fa1889(ip_38_26,ip_39_25,ip_40_24,p5910,p5911);
FA fa1890(ip_41_23,ip_42_22,ip_43_21,p5912,p5913);
HA ha1066(ip_44_20,ip_45_19,p5914,p5915);
FA fa1891(ip_46_18,ip_47_17,ip_48_16,p5916,p5917);
HA ha1067(ip_49_15,ip_50_14,p5918,p5919);
FA fa1892(ip_51_13,ip_52_12,ip_53_11,p5920,p5921);
FA fa1893(ip_54_10,ip_55_9,ip_56_8,p5922,p5923);
FA fa1894(ip_57_7,ip_58_6,ip_59_5,p5924,p5925);
FA fa1895(ip_60_4,ip_61_3,ip_62_2,p5926,p5927);
HA ha1068(ip_63_1,p5694,p5928,p5929);
HA ha1069(p5708,p5714,p5930,p5931);
FA fa1896(p5720,p5728,p5732,p5932,p5933);
FA fa1897(p5734,p5887,p5889,p5934,p5935);
FA fa1898(p5891,p5901,p5905,p5936,p5937);
FA fa1899(p5915,p5919,p5740,p5938,p5939);
FA fa1900(p5746,p5748,p5883,p5940,p5941);
FA fa1901(p5885,p5893,p5895,p5942,p5943);
HA ha1070(p5897,p5899,p5944,p5945);
FA fa1902(p5903,p5907,p5909,p5946,p5947);
HA ha1071(p5911,p5913,p5948,p5949);
HA ha1072(p5917,p5921,p5950,p5951);
FA fa1903(p5923,p5925,p5927,p5952,p5953);
FA fa1904(p5929,p5931,p5690,p5954,p5955);
HA ha1073(p5692,p5696,p5956,p5957);
FA fa1905(p5698,p5700,p5702,p5958,p5959);
HA ha1074(p5704,p5706,p5960,p5961);
HA ha1075(p5710,p5712,p5962,p5963);
FA fa1906(p5716,p5718,p5722,p5964,p5965);
FA fa1907(p5724,p5726,p5730,p5966,p5967);
FA fa1908(p5736,p5750,p5756,p5968,p5969);
FA fa1909(p5764,p5933,p5935,p5970,p5971);
HA ha1076(p5937,p5939,p5972,p5973);
FA fa1910(p5945,p5949,p5951,p5974,p5975);
HA ha1077(p5738,p5742,p5976,p5977);
FA fa1911(p5744,p5782,p5941,p5978,p5979);
FA fa1912(p5943,p5947,p5953,p5980,p5981);
FA fa1913(p5955,p5957,p5961,p5982,p5983);
FA fa1914(p5963,p5973,p5752,p5984,p5985);
FA fa1915(p5754,p5758,p5760,p5986,p5987);
HA ha1078(p5762,p5766,p5988,p5989);
FA fa1916(p5784,p5788,p5790,p5990,p5991);
FA fa1917(p5959,p5965,p5967,p5992,p5993);
FA fa1918(p5969,p5971,p5975,p5994,p5995);
FA fa1919(p5977,p5768,p5770,p5996,p5997);
FA fa1920(p5772,p5774,p5776,p5998,p5999);
FA fa1921(p5778,p5780,p5798,p6000,p6001);
FA fa1922(p5802,p5979,p5981,p6002,p6003);
FA fa1923(p5983,p5985,p5989,p6004,p6005);
HA ha1079(p5786,p5792,p6006,p6007);
FA fa1924(p5794,p5987,p5991,p6008,p6009);
FA fa1925(p5993,p5995,p5796,p6010,p6011);
HA ha1080(p5800,p5804,p6012,p6013);
HA ha1081(p5806,p5997,p6014,p6015);
FA fa1926(p5999,p6001,p6003,p6016,p6017);
FA fa1927(p6005,p6007,p5808,p6018,p6019);
HA ha1082(p5810,p5812,p6020,p6021);
HA ha1083(p5814,p5822,p6022,p6023);
HA ha1084(p5828,p6009,p6024,p6025);
HA ha1085(p6011,p6013,p6026,p6027);
FA fa1928(p6015,p5816,p5818,p6028,p6029);
HA ha1086(p5834,p5838,p6030,p6031);
FA fa1929(p6017,p6019,p6021,p6032,p6033);
FA fa1930(p6023,p6025,p6027,p6034,p6035);
HA ha1087(p5820,p5824,p6036,p6037);
FA fa1931(p5826,p5840,p5846,p6038,p6039);
FA fa1932(p6031,p5830,p5832,p6040,p6041);
HA ha1088(p5836,p6029,p6042,p6043);
HA ha1089(p6033,p6035,p6044,p6045);
HA ha1090(p6037,p5842,p6046,p6047);
FA fa1933(p5844,p6039,p6043,p6048,p6049);
FA fa1934(p6045,p5848,p5850,p6050,p6051);
HA ha1091(p5858,p6041,p6052,p6053);
FA fa1935(p6047,p5852,p5854,p6054,p6055);
FA fa1936(p5864,p6049,p6053,p6056,p6057);
HA ha1092(p5856,p6051,p6058,p6059);
FA fa1937(p5860,p5862,p6055,p6060,p6061);
FA fa1938(p6057,p6059,p5866,p6062,p6063);
HA ha1093(p5870,p5872,p6064,p6065);
FA fa1939(p5868,p6061,p6063,p6066,p6067);
FA fa1940(p6065,p5874,p6067,p6068,p6069);
HA ha1094(p5876,p6069,p6070,p6071);
FA fa1941(p5878,p6071,p5880,p6072,p6073);
FA fa1942(ip_2_63,ip_3_62,ip_4_61,p6074,p6075);
FA fa1943(ip_5_60,ip_6_59,ip_7_58,p6076,p6077);
FA fa1944(ip_8_57,ip_9_56,ip_10_55,p6078,p6079);
FA fa1945(ip_11_54,ip_12_53,ip_13_52,p6080,p6081);
HA ha1095(ip_14_51,ip_15_50,p6082,p6083);
FA fa1946(ip_16_49,ip_17_48,ip_18_47,p6084,p6085);
FA fa1947(ip_19_46,ip_20_45,ip_21_44,p6086,p6087);
FA fa1948(ip_22_43,ip_23_42,ip_24_41,p6088,p6089);
FA fa1949(ip_25_40,ip_26_39,ip_27_38,p6090,p6091);
HA ha1096(ip_28_37,ip_29_36,p6092,p6093);
FA fa1950(ip_30_35,ip_31_34,ip_32_33,p6094,p6095);
HA ha1097(ip_33_32,ip_34_31,p6096,p6097);
FA fa1951(ip_35_30,ip_36_29,ip_37_28,p6098,p6099);
FA fa1952(ip_38_27,ip_39_26,ip_40_25,p6100,p6101);
HA ha1098(ip_41_24,ip_42_23,p6102,p6103);
FA fa1953(ip_43_22,ip_44_21,ip_45_20,p6104,p6105);
HA ha1099(ip_46_19,ip_47_18,p6106,p6107);
FA fa1954(ip_48_17,ip_49_16,ip_50_15,p6108,p6109);
FA fa1955(ip_51_14,ip_52_13,ip_53_12,p6110,p6111);
FA fa1956(ip_54_11,ip_55_10,ip_56_9,p6112,p6113);
FA fa1957(ip_57_8,ip_58_7,ip_59_6,p6114,p6115);
FA fa1958(ip_60_5,ip_61_4,ip_62_3,p6116,p6117);
HA ha1100(ip_63_2,p5886,p6118,p6119);
FA fa1959(p5888,p5890,p5900,p6120,p6121);
FA fa1960(p5904,p5914,p5918,p6122,p6123);
HA ha1101(p6083,p6093,p6124,p6125);
HA ha1102(p6097,p6103,p6126,p6127);
HA ha1103(p6107,p5928,p6128,p6129);
HA ha1104(p5930,p6075,p6130,p6131);
FA fa1961(p6077,p6079,p6081,p6132,p6133);
FA fa1962(p6085,p6087,p6089,p6134,p6135);
FA fa1963(p6091,p6095,p6099,p6136,p6137);
FA fa1964(p6101,p6105,p6109,p6138,p6139);
FA fa1965(p6111,p6113,p6115,p6140,p6141);
FA fa1966(p6117,p6119,p6125,p6142,p6143);
FA fa1967(p6127,p5882,p5884,p6144,p6145);
HA ha1105(p5892,p5894,p6146,p6147);
FA fa1968(p5896,p5898,p5902,p6148,p6149);
FA fa1969(p5906,p5908,p5910,p6150,p6151);
FA fa1970(p5912,p5916,p5920,p6152,p6153);
HA ha1106(p5922,p5924,p6154,p6155);
FA fa1971(p5926,p5944,p5948,p6156,p6157);
FA fa1972(p5950,p6121,p6123,p6158,p6159);
HA ha1107(p6129,p6131,p6160,p6161);
FA fa1973(p5932,p5934,p5936,p6162,p6163);
FA fa1974(p5938,p5956,p5960,p6164,p6165);
FA fa1975(p5962,p5972,p6133,p6166,p6167);
HA ha1108(p6135,p6137,p6168,p6169);
HA ha1109(p6139,p6141,p6170,p6171);
FA fa1976(p6143,p6147,p6155,p6172,p6173);
FA fa1977(p6161,p5940,p5942,p6174,p6175);
FA fa1978(p5946,p5952,p5954,p6176,p6177);
HA ha1110(p5976,p6145,p6178,p6179);
HA ha1111(p6149,p6151,p6180,p6181);
FA fa1979(p6153,p6157,p6159,p6182,p6183);
FA fa1980(p6169,p6171,p5958,p6184,p6185);
FA fa1981(p5964,p5966,p5968,p6186,p6187);
FA fa1982(p5970,p5974,p5988,p6188,p6189);
FA fa1983(p6163,p6165,p6167,p6190,p6191);
FA fa1984(p6173,p6179,p6181,p6192,p6193);
FA fa1985(p5978,p5980,p5982,p6194,p6195);
FA fa1986(p5984,p6175,p6177,p6196,p6197);
FA fa1987(p6183,p6185,p5986,p6198,p6199);
FA fa1988(p5990,p5992,p5994,p6200,p6201);
FA fa1989(p6006,p6187,p6189,p6202,p6203);
HA ha1112(p6191,p6193,p6204,p6205);
FA fa1990(p5996,p5998,p6000,p6206,p6207);
FA fa1991(p6002,p6004,p6012,p6208,p6209);
FA fa1992(p6014,p6195,p6197,p6210,p6211);
HA ha1113(p6199,p6205,p6212,p6213);
HA ha1114(p6008,p6010,p6214,p6215);
FA fa1993(p6020,p6022,p6024,p6216,p6217);
FA fa1994(p6026,p6201,p6203,p6218,p6219);
FA fa1995(p6213,p6016,p6018,p6220,p6221);
FA fa1996(p6030,p6207,p6209,p6222,p6223);
HA ha1115(p6211,p6215,p6224,p6225);
FA fa1997(p6036,p6217,p6219,p6226,p6227);
HA ha1116(p6225,p6028,p6228,p6229);
FA fa1998(p6032,p6034,p6042,p6230,p6231);
FA fa1999(p6044,p6221,p6223,p6232,p6233);
HA ha1117(p6038,p6046,p6234,p6235);
FA fa2000(p6227,p6229,p6040,p6236,p6237);
FA fa2001(p6052,p6231,p6233,p6238,p6239);
HA ha1118(p6235,p6048,p6240,p6241);
HA ha1119(p6237,p6050,p6242,p6243);
HA ha1120(p6058,p6239,p6244,p6245);
FA fa2002(p6241,p6054,p6056,p6246,p6247);
HA ha1121(p6243,p6245,p6248,p6249);
FA fa2003(p6064,p6249,p6060,p6250,p6251);
FA fa2004(p6062,p6247,p6251,p6252,p6253);
FA fa2005(p6066,p6253,p6068,p6254,p6255);
FA fa2006(p6070,p6255,p6072,p6256,p6257);
HA ha1122(ip_3_63,ip_4_62,p6258,p6259);
FA fa2007(ip_5_61,ip_6_60,ip_7_59,p6260,p6261);
FA fa2008(ip_8_58,ip_9_57,ip_10_56,p6262,p6263);
FA fa2009(ip_11_55,ip_12_54,ip_13_53,p6264,p6265);
FA fa2010(ip_14_52,ip_15_51,ip_16_50,p6266,p6267);
FA fa2011(ip_17_49,ip_18_48,ip_19_47,p6268,p6269);
FA fa2012(ip_20_46,ip_21_45,ip_22_44,p6270,p6271);
FA fa2013(ip_23_43,ip_24_42,ip_25_41,p6272,p6273);
FA fa2014(ip_26_40,ip_27_39,ip_28_38,p6274,p6275);
HA ha1123(ip_29_37,ip_30_36,p6276,p6277);
FA fa2015(ip_31_35,ip_32_34,ip_33_33,p6278,p6279);
FA fa2016(ip_34_32,ip_35_31,ip_36_30,p6280,p6281);
FA fa2017(ip_37_29,ip_38_28,ip_39_27,p6282,p6283);
FA fa2018(ip_40_26,ip_41_25,ip_42_24,p6284,p6285);
FA fa2019(ip_43_23,ip_44_22,ip_45_21,p6286,p6287);
HA ha1124(ip_46_20,ip_47_19,p6288,p6289);
HA ha1125(ip_48_18,ip_49_17,p6290,p6291);
FA fa2020(ip_50_16,ip_51_15,ip_52_14,p6292,p6293);
FA fa2021(ip_53_13,ip_54_12,ip_55_11,p6294,p6295);
FA fa2022(ip_56_10,ip_57_9,ip_58_8,p6296,p6297);
HA ha1126(ip_59_7,ip_60_6,p6298,p6299);
HA ha1127(ip_61_5,ip_62_4,p6300,p6301);
FA fa2023(ip_63_3,p6082,p6092,p6302,p6303);
FA fa2024(p6096,p6102,p6106,p6304,p6305);
FA fa2025(p6259,p6277,p6289,p6306,p6307);
HA ha1128(p6291,p6299,p6308,p6309);
HA ha1129(p6301,p6118,p6310,p6311);
FA fa2026(p6124,p6126,p6261,p6312,p6313);
FA fa2027(p6263,p6265,p6267,p6314,p6315);
HA ha1130(p6269,p6271,p6316,p6317);
HA ha1131(p6273,p6275,p6318,p6319);
FA fa2028(p6279,p6281,p6283,p6320,p6321);
FA fa2029(p6285,p6287,p6293,p6322,p6323);
FA fa2030(p6295,p6297,p6309,p6324,p6325);
FA fa2031(p6074,p6076,p6078,p6326,p6327);
FA fa2032(p6080,p6084,p6086,p6328,p6329);
HA ha1132(p6088,p6090,p6330,p6331);
HA ha1133(p6094,p6098,p6332,p6333);
FA fa2033(p6100,p6104,p6108,p6334,p6335);
HA ha1134(p6110,p6112,p6336,p6337);
HA ha1135(p6114,p6116,p6338,p6339);
FA fa2034(p6128,p6130,p6303,p6340,p6341);
FA fa2035(p6305,p6307,p6311,p6342,p6343);
FA fa2036(p6317,p6319,p6120,p6344,p6345);
HA ha1136(p6122,p6146,p6346,p6347);
FA fa2037(p6154,p6160,p6313,p6348,p6349);
HA ha1137(p6315,p6321,p6350,p6351);
FA fa2038(p6323,p6325,p6331,p6352,p6353);
FA fa2039(p6333,p6337,p6339,p6354,p6355);
FA fa2040(p6132,p6134,p6136,p6356,p6357);
HA ha1138(p6138,p6140,p6358,p6359);
FA fa2041(p6142,p6168,p6170,p6360,p6361);
FA fa2042(p6327,p6329,p6335,p6362,p6363);
HA ha1139(p6341,p6343,p6364,p6365);
FA fa2043(p6345,p6347,p6351,p6366,p6367);
FA fa2044(p6144,p6148,p6150,p6368,p6369);
HA ha1140(p6152,p6156,p6370,p6371);
FA fa2045(p6158,p6178,p6180,p6372,p6373);
FA fa2046(p6349,p6353,p6355,p6374,p6375);
FA fa2047(p6359,p6365,p6162,p6376,p6377);
FA fa2048(p6164,p6166,p6172,p6378,p6379);
FA fa2049(p6357,p6361,p6363,p6380,p6381);
FA fa2050(p6367,p6371,p6174,p6382,p6383);
HA ha1141(p6176,p6182,p6384,p6385);
FA fa2051(p6184,p6369,p6373,p6386,p6387);
FA fa2052(p6375,p6377,p6186,p6388,p6389);
FA fa2053(p6188,p6190,p6192,p6390,p6391);
FA fa2054(p6204,p6379,p6381,p6392,p6393);
HA ha1142(p6383,p6385,p6394,p6395);
HA ha1143(p6194,p6196,p6396,p6397);
HA ha1144(p6198,p6212,p6398,p6399);
FA fa2055(p6387,p6389,p6395,p6400,p6401);
HA ha1145(p6200,p6202,p6402,p6403);
FA fa2056(p6214,p6391,p6393,p6404,p6405);
HA ha1146(p6397,p6399,p6406,p6407);
HA ha1147(p6206,p6208,p6408,p6409);
HA ha1148(p6210,p6224,p6410,p6411);
HA ha1149(p6401,p6403,p6412,p6413);
HA ha1150(p6407,p6216,p6414,p6415);
FA fa2057(p6218,p6405,p6409,p6416,p6417);
FA fa2058(p6411,p6413,p6220,p6418,p6419);
FA fa2059(p6222,p6228,p6415,p6420,p6421);
FA fa2060(p6226,p6234,p6417,p6422,p6423);
FA fa2061(p6419,p6230,p6232,p6424,p6425);
HA ha1151(p6421,p6236,p6426,p6427);
FA fa2062(p6240,p6423,p6238,p6428,p6429);
FA fa2063(p6242,p6244,p6425,p6430,p6431);
FA fa2064(p6427,p6248,p6429,p6432,p6433);
HA ha1152(p6431,p6246,p6434,p6435);
HA ha1153(p6433,p6250,p6436,p6437);
FA fa2065(p6435,p6252,p6437,p6438,p6439);
FA fa2066(p6439,p6254,p6256,p6440,p6441);
HA ha1154(ip_4_63,ip_5_62,p6442,p6443);
FA fa2067(ip_6_61,ip_7_60,ip_8_59,p6444,p6445);
FA fa2068(ip_9_58,ip_10_57,ip_11_56,p6446,p6447);
FA fa2069(ip_12_55,ip_13_54,ip_14_53,p6448,p6449);
FA fa2070(ip_15_52,ip_16_51,ip_17_50,p6450,p6451);
HA ha1155(ip_18_49,ip_19_48,p6452,p6453);
HA ha1156(ip_20_47,ip_21_46,p6454,p6455);
FA fa2071(ip_22_45,ip_23_44,ip_24_43,p6456,p6457);
HA ha1157(ip_25_42,ip_26_41,p6458,p6459);
FA fa2072(ip_27_40,ip_28_39,ip_29_38,p6460,p6461);
FA fa2073(ip_30_37,ip_31_36,ip_32_35,p6462,p6463);
HA ha1158(ip_33_34,ip_34_33,p6464,p6465);
HA ha1159(ip_35_32,ip_36_31,p6466,p6467);
HA ha1160(ip_37_30,ip_38_29,p6468,p6469);
FA fa2074(ip_39_28,ip_40_27,ip_41_26,p6470,p6471);
FA fa2075(ip_42_25,ip_43_24,ip_44_23,p6472,p6473);
FA fa2076(ip_45_22,ip_46_21,ip_47_20,p6474,p6475);
HA ha1161(ip_48_19,ip_49_18,p6476,p6477);
HA ha1162(ip_50_17,ip_51_16,p6478,p6479);
FA fa2077(ip_52_15,ip_53_14,ip_54_13,p6480,p6481);
HA ha1163(ip_55_12,ip_56_11,p6482,p6483);
FA fa2078(ip_57_10,ip_58_9,ip_59_8,p6484,p6485);
FA fa2079(ip_60_7,ip_61_6,ip_62_5,p6486,p6487);
FA fa2080(ip_63_4,p6258,p6276,p6488,p6489);
FA fa2081(p6288,p6290,p6298,p6490,p6491);
HA ha1164(p6300,p6443,p6492,p6493);
FA fa2082(p6453,p6455,p6459,p6494,p6495);
FA fa2083(p6465,p6467,p6469,p6496,p6497);
FA fa2084(p6477,p6479,p6483,p6498,p6499);
HA ha1165(p6308,p6445,p6500,p6501);
HA ha1166(p6447,p6449,p6502,p6503);
HA ha1167(p6451,p6457,p6504,p6505);
FA fa2085(p6461,p6463,p6471,p6506,p6507);
FA fa2086(p6473,p6475,p6481,p6508,p6509);
FA fa2087(p6485,p6487,p6493,p6510,p6511);
HA ha1168(p6260,p6262,p6512,p6513);
HA ha1169(p6264,p6266,p6514,p6515);
FA fa2088(p6268,p6270,p6272,p6516,p6517);
FA fa2089(p6274,p6278,p6280,p6518,p6519);
HA ha1170(p6282,p6284,p6520,p6521);
FA fa2090(p6286,p6292,p6294,p6522,p6523);
FA fa2091(p6296,p6310,p6316,p6524,p6525);
HA ha1171(p6318,p6489,p6526,p6527);
HA ha1172(p6491,p6495,p6528,p6529);
HA ha1173(p6497,p6499,p6530,p6531);
FA fa2092(p6501,p6503,p6505,p6532,p6533);
FA fa2093(p6302,p6304,p6306,p6534,p6535);
FA fa2094(p6330,p6332,p6336,p6536,p6537);
FA fa2095(p6338,p6507,p6509,p6538,p6539);
FA fa2096(p6511,p6513,p6515,p6540,p6541);
FA fa2097(p6521,p6527,p6529,p6542,p6543);
HA ha1174(p6531,p6312,p6544,p6545);
FA fa2098(p6314,p6320,p6322,p6546,p6547);
FA fa2099(p6324,p6346,p6350,p6548,p6549);
FA fa2100(p6517,p6519,p6523,p6550,p6551);
FA fa2101(p6525,p6533,p6326,p6552,p6553);
HA ha1175(p6328,p6334,p6554,p6555);
HA ha1176(p6340,p6342,p6556,p6557);
FA fa2102(p6344,p6358,p6364,p6558,p6559);
FA fa2103(p6535,p6537,p6539,p6560,p6561);
HA ha1177(p6541,p6543,p6562,p6563);
HA ha1178(p6545,p6348,p6564,p6565);
FA fa2104(p6352,p6354,p6370,p6566,p6567);
HA ha1179(p6547,p6549,p6568,p6569);
FA fa2105(p6551,p6553,p6555,p6570,p6571);
FA fa2106(p6557,p6563,p6356,p6572,p6573);
FA fa2107(p6360,p6362,p6366,p6574,p6575);
FA fa2108(p6559,p6561,p6565,p6576,p6577);
FA fa2109(p6569,p6368,p6372,p6578,p6579);
FA fa2110(p6374,p6376,p6384,p6580,p6581);
FA fa2111(p6567,p6571,p6573,p6582,p6583);
HA ha1180(p6378,p6380,p6584,p6585);
FA fa2112(p6382,p6394,p6575,p6586,p6587);
FA fa2113(p6577,p6386,p6388,p6588,p6589);
FA fa2114(p6396,p6398,p6579,p6590,p6591);
FA fa2115(p6581,p6583,p6585,p6592,p6593);
FA fa2116(p6390,p6392,p6402,p6594,p6595);
FA fa2117(p6406,p6587,p6400,p6596,p6597);
HA ha1181(p6408,p6410,p6598,p6599);
HA ha1182(p6412,p6589,p6600,p6601);
FA fa2118(p6591,p6593,p6404,p6602,p6603);
FA fa2119(p6414,p6595,p6597,p6604,p6605);
HA ha1183(p6599,p6601,p6606,p6607);
FA fa2120(p6603,p6607,p6416,p6608,p6609);
FA fa2121(p6418,p6605,p6420,p6610,p6611);
FA fa2122(p6609,p6422,p6426,p6612,p6613);
HA ha1184(p6611,p6424,p6614,p6615);
FA fa2123(p6428,p6613,p6615,p6616,p6617);
HA ha1185(p6430,p6432,p6618,p6619);
FA fa2124(p6434,p6617,p6436,p6620,p6621);
FA fa2125(p6619,p6621,p6438,p6622,p6623);
HA ha1186(ip_5_63,ip_6_62,p6624,p6625);
HA ha1187(ip_7_61,ip_8_60,p6626,p6627);
FA fa2126(ip_9_59,ip_10_58,ip_11_57,p6628,p6629);
HA ha1188(ip_12_56,ip_13_55,p6630,p6631);
FA fa2127(ip_14_54,ip_15_53,ip_16_52,p6632,p6633);
FA fa2128(ip_17_51,ip_18_50,ip_19_49,p6634,p6635);
FA fa2129(ip_20_48,ip_21_47,ip_22_46,p6636,p6637);
FA fa2130(ip_23_45,ip_24_44,ip_25_43,p6638,p6639);
FA fa2131(ip_26_42,ip_27_41,ip_28_40,p6640,p6641);
FA fa2132(ip_29_39,ip_30_38,ip_31_37,p6642,p6643);
FA fa2133(ip_32_36,ip_33_35,ip_34_34,p6644,p6645);
HA ha1189(ip_35_33,ip_36_32,p6646,p6647);
HA ha1190(ip_37_31,ip_38_30,p6648,p6649);
HA ha1191(ip_39_29,ip_40_28,p6650,p6651);
FA fa2134(ip_41_27,ip_42_26,ip_43_25,p6652,p6653);
FA fa2135(ip_44_24,ip_45_23,ip_46_22,p6654,p6655);
HA ha1192(ip_47_21,ip_48_20,p6656,p6657);
HA ha1193(ip_49_19,ip_50_18,p6658,p6659);
FA fa2136(ip_51_17,ip_52_16,ip_53_15,p6660,p6661);
HA ha1194(ip_54_14,ip_55_13,p6662,p6663);
FA fa2137(ip_56_12,ip_57_11,ip_58_10,p6664,p6665);
HA ha1195(ip_59_9,ip_60_8,p6666,p6667);
FA fa2138(ip_61_7,ip_62_6,ip_63_5,p6668,p6669);
FA fa2139(p6442,p6452,p6454,p6670,p6671);
FA fa2140(p6458,p6464,p6466,p6672,p6673);
FA fa2141(p6468,p6476,p6478,p6674,p6675);
FA fa2142(p6482,p6625,p6627,p6676,p6677);
FA fa2143(p6631,p6647,p6649,p6678,p6679);
FA fa2144(p6651,p6657,p6659,p6680,p6681);
HA ha1196(p6663,p6667,p6682,p6683);
HA ha1197(p6492,p6629,p6684,p6685);
FA fa2145(p6633,p6635,p6637,p6686,p6687);
FA fa2146(p6639,p6641,p6643,p6688,p6689);
FA fa2147(p6645,p6653,p6655,p6690,p6691);
HA ha1198(p6661,p6665,p6692,p6693);
HA ha1199(p6669,p6683,p6694,p6695);
FA fa2148(p6444,p6446,p6448,p6696,p6697);
FA fa2149(p6450,p6456,p6460,p6698,p6699);
FA fa2150(p6462,p6470,p6472,p6700,p6701);
HA ha1200(p6474,p6480,p6702,p6703);
FA fa2151(p6484,p6486,p6500,p6704,p6705);
FA fa2152(p6502,p6504,p6671,p6706,p6707);
FA fa2153(p6673,p6675,p6677,p6708,p6709);
HA ha1201(p6679,p6681,p6710,p6711);
FA fa2154(p6685,p6693,p6695,p6712,p6713);
FA fa2155(p6488,p6490,p6494,p6714,p6715);
HA ha1202(p6496,p6498,p6716,p6717);
FA fa2156(p6512,p6514,p6520,p6718,p6719);
HA ha1203(p6526,p6528,p6720,p6721);
HA ha1204(p6530,p6687,p6722,p6723);
HA ha1205(p6689,p6691,p6724,p6725);
FA fa2157(p6703,p6711,p6506,p6726,p6727);
HA ha1206(p6508,p6510,p6728,p6729);
FA fa2158(p6697,p6699,p6701,p6730,p6731);
FA fa2159(p6705,p6707,p6709,p6732,p6733);
FA fa2160(p6713,p6717,p6721,p6734,p6735);
FA fa2161(p6723,p6725,p6516,p6736,p6737);
FA fa2162(p6518,p6522,p6524,p6738,p6739);
FA fa2163(p6532,p6544,p6715,p6740,p6741);
HA ha1207(p6719,p6727,p6742,p6743);
FA fa2164(p6729,p6534,p6536,p6744,p6745);
FA fa2165(p6538,p6540,p6542,p6746,p6747);
FA fa2166(p6554,p6556,p6562,p6748,p6749);
FA fa2167(p6731,p6733,p6735,p6750,p6751);
HA ha1208(p6737,p6743,p6752,p6753);
FA fa2168(p6546,p6548,p6550,p6754,p6755);
FA fa2169(p6552,p6564,p6568,p6756,p6757);
HA ha1209(p6739,p6741,p6758,p6759);
HA ha1210(p6753,p6558,p6760,p6761);
HA ha1211(p6560,p6745,p6762,p6763);
FA fa2170(p6747,p6749,p6751,p6764,p6765);
HA ha1212(p6759,p6566,p6766,p6767);
HA ha1213(p6570,p6572,p6768,p6769);
FA fa2171(p6755,p6757,p6761,p6770,p6771);
FA fa2172(p6763,p6574,p6576,p6772,p6773);
HA ha1214(p6584,p6765,p6774,p6775);
HA ha1215(p6767,p6769,p6776,p6777);
HA ha1216(p6578,p6580,p6778,p6779);
FA fa2173(p6582,p6771,p6775,p6780,p6781);
FA fa2174(p6777,p6586,p6773,p6782,p6783);
FA fa2175(p6779,p6588,p6590,p6784,p6785);
FA fa2176(p6592,p6598,p6600,p6786,p6787);
FA fa2177(p6781,p6594,p6596,p6788,p6789);
FA fa2178(p6606,p6783,p6602,p6790,p6791);
HA ha1217(p6785,p6787,p6792,p6793);
HA ha1218(p6604,p6789,p6794,p6795);
FA fa2179(p6791,p6793,p6608,p6796,p6797);
FA fa2180(p6795,p6610,p6797,p6798,p6799);
HA ha1219(p6614,p6612,p6800,p6801);
HA ha1220(p6799,p6801,p6802,p6803);
FA fa2181(p6616,p6618,p6803,p6804,p6805);
FA fa2182(p6620,p6805,p6622,p6806,p6807);
FA fa2183(ip_6_63,ip_7_62,ip_8_61,p6808,p6809);
FA fa2184(ip_9_60,ip_10_59,ip_11_58,p6810,p6811);
FA fa2185(ip_12_57,ip_13_56,ip_14_55,p6812,p6813);
HA ha1221(ip_15_54,ip_16_53,p6814,p6815);
FA fa2186(ip_17_52,ip_18_51,ip_19_50,p6816,p6817);
HA ha1222(ip_20_49,ip_21_48,p6818,p6819);
FA fa2187(ip_22_47,ip_23_46,ip_24_45,p6820,p6821);
FA fa2188(ip_25_44,ip_26_43,ip_27_42,p6822,p6823);
HA ha1223(ip_28_41,ip_29_40,p6824,p6825);
FA fa2189(ip_30_39,ip_31_38,ip_32_37,p6826,p6827);
FA fa2190(ip_33_36,ip_34_35,ip_35_34,p6828,p6829);
FA fa2191(ip_36_33,ip_37_32,ip_38_31,p6830,p6831);
HA ha1224(ip_39_30,ip_40_29,p6832,p6833);
FA fa2192(ip_41_28,ip_42_27,ip_43_26,p6834,p6835);
FA fa2193(ip_44_25,ip_45_24,ip_46_23,p6836,p6837);
FA fa2194(ip_47_22,ip_48_21,ip_49_20,p6838,p6839);
FA fa2195(ip_50_19,ip_51_18,ip_52_17,p6840,p6841);
FA fa2196(ip_53_16,ip_54_15,ip_55_14,p6842,p6843);
FA fa2197(ip_56_13,ip_57_12,ip_58_11,p6844,p6845);
FA fa2198(ip_59_10,ip_60_9,ip_61_8,p6846,p6847);
FA fa2199(ip_62_7,ip_63_6,p6624,p6848,p6849);
HA ha1225(p6626,p6630,p6850,p6851);
FA fa2200(p6646,p6648,p6650,p6852,p6853);
FA fa2201(p6656,p6658,p6662,p6854,p6855);
FA fa2202(p6666,p6815,p6819,p6856,p6857);
HA ha1226(p6825,p6833,p6858,p6859);
FA fa2203(p6682,p6809,p6811,p6860,p6861);
HA ha1227(p6813,p6817,p6862,p6863);
HA ha1228(p6821,p6823,p6864,p6865);
FA fa2204(p6827,p6829,p6831,p6866,p6867);
HA ha1229(p6835,p6837,p6868,p6869);
FA fa2205(p6839,p6841,p6843,p6870,p6871);
FA fa2206(p6845,p6847,p6849,p6872,p6873);
FA fa2207(p6851,p6859,p6628,p6874,p6875);
FA fa2208(p6632,p6634,p6636,p6876,p6877);
HA ha1230(p6638,p6640,p6878,p6879);
HA ha1231(p6642,p6644,p6880,p6881);
FA fa2209(p6652,p6654,p6660,p6882,p6883);
HA ha1232(p6664,p6668,p6884,p6885);
FA fa2210(p6684,p6692,p6694,p6886,p6887);
FA fa2211(p6853,p6855,p6857,p6888,p6889);
FA fa2212(p6863,p6865,p6869,p6890,p6891);
FA fa2213(p6670,p6672,p6674,p6892,p6893);
FA fa2214(p6676,p6678,p6680,p6894,p6895);
FA fa2215(p6702,p6710,p6861,p6896,p6897);
FA fa2216(p6867,p6871,p6873,p6898,p6899);
FA fa2217(p6875,p6879,p6881,p6900,p6901);
HA ha1233(p6885,p6686,p6902,p6903);
FA fa2218(p6688,p6690,p6716,p6904,p6905);
FA fa2219(p6720,p6722,p6724,p6906,p6907);
HA ha1234(p6877,p6883,p6908,p6909);
HA ha1235(p6887,p6889,p6910,p6911);
FA fa2220(p6891,p6696,p6698,p6912,p6913);
FA fa2221(p6700,p6704,p6706,p6914,p6915);
FA fa2222(p6708,p6712,p6728,p6916,p6917);
FA fa2223(p6893,p6895,p6897,p6918,p6919);
FA fa2224(p6899,p6901,p6903,p6920,p6921);
FA fa2225(p6909,p6911,p6714,p6922,p6923);
FA fa2226(p6718,p6726,p6742,p6924,p6925);
FA fa2227(p6905,p6907,p6730,p6926,p6927);
HA ha1236(p6732,p6734,p6928,p6929);
HA ha1237(p6736,p6752,p6930,p6931);
FA fa2228(p6913,p6915,p6917,p6932,p6933);
FA fa2229(p6919,p6921,p6923,p6934,p6935);
FA fa2230(p6738,p6740,p6758,p6936,p6937);
HA ha1238(p6925,p6927,p6938,p6939);
FA fa2231(p6929,p6931,p6744,p6940,p6941);
FA fa2232(p6746,p6748,p6750,p6942,p6943);
FA fa2233(p6760,p6762,p6933,p6944,p6945);
FA fa2234(p6935,p6939,p6754,p6946,p6947);
HA ha1239(p6756,p6766,p6948,p6949);
FA fa2235(p6768,p6937,p6941,p6950,p6951);
FA fa2236(p6764,p6774,p6776,p6952,p6953);
FA fa2237(p6943,p6945,p6947,p6954,p6955);
HA ha1240(p6949,p6770,p6956,p6957);
HA ha1241(p6778,p6951,p6958,p6959);
FA fa2238(p6772,p6953,p6955,p6960,p6961);
FA fa2239(p6957,p6959,p6780,p6962,p6963);
HA ha1242(p6782,p6961,p6964,p6965);
FA fa2240(p6963,p6784,p6786,p6966,p6967);
FA fa2241(p6792,p6965,p6788,p6968,p6969);
FA fa2242(p6790,p6794,p6967,p6970,p6971);
FA fa2243(p6969,p6796,p6971,p6972,p6973);
FA fa2244(p6798,p6800,p6973,p6974,p6975);
FA fa2245(p6802,p6975,p6804,p6976,p6977);
HA ha1243(ip_7_63,ip_8_62,p6978,p6979);
FA fa2246(ip_9_61,ip_10_60,ip_11_59,p6980,p6981);
FA fa2247(ip_12_58,ip_13_57,ip_14_56,p6982,p6983);
HA ha1244(ip_15_55,ip_16_54,p6984,p6985);
FA fa2248(ip_17_53,ip_18_52,ip_19_51,p6986,p6987);
HA ha1245(ip_20_50,ip_21_49,p6988,p6989);
FA fa2249(ip_22_48,ip_23_47,ip_24_46,p6990,p6991);
FA fa2250(ip_25_45,ip_26_44,ip_27_43,p6992,p6993);
HA ha1246(ip_28_42,ip_29_41,p6994,p6995);
FA fa2251(ip_30_40,ip_31_39,ip_32_38,p6996,p6997);
HA ha1247(ip_33_37,ip_34_36,p6998,p6999);
HA ha1248(ip_35_35,ip_36_34,p7000,p7001);
FA fa2252(ip_37_33,ip_38_32,ip_39_31,p7002,p7003);
FA fa2253(ip_40_30,ip_41_29,ip_42_28,p7004,p7005);
FA fa2254(ip_43_27,ip_44_26,ip_45_25,p7006,p7007);
FA fa2255(ip_46_24,ip_47_23,ip_48_22,p7008,p7009);
FA fa2256(ip_49_21,ip_50_20,ip_51_19,p7010,p7011);
HA ha1249(ip_52_18,ip_53_17,p7012,p7013);
HA ha1250(ip_54_16,ip_55_15,p7014,p7015);
FA fa2257(ip_56_14,ip_57_13,ip_58_12,p7016,p7017);
FA fa2258(ip_59_11,ip_60_10,ip_61_9,p7018,p7019);
FA fa2259(ip_62_8,ip_63_7,p6814,p7020,p7021);
FA fa2260(p6818,p6824,p6832,p7022,p7023);
FA fa2261(p6979,p6985,p6989,p7024,p7025);
FA fa2262(p6995,p6999,p7001,p7026,p7027);
HA ha1251(p7013,p7015,p7028,p7029);
FA fa2263(p6850,p6858,p6981,p7030,p7031);
FA fa2264(p6983,p6987,p6991,p7032,p7033);
HA ha1252(p6993,p6997,p7034,p7035);
FA fa2265(p7003,p7005,p7007,p7036,p7037);
FA fa2266(p7009,p7011,p7017,p7038,p7039);
HA ha1253(p7019,p7021,p7040,p7041);
FA fa2267(p7029,p6808,p6810,p7042,p7043);
FA fa2268(p6812,p6816,p6820,p7044,p7045);
FA fa2269(p6822,p6826,p6828,p7046,p7047);
FA fa2270(p6830,p6834,p6836,p7048,p7049);
HA ha1254(p6838,p6840,p7050,p7051);
HA ha1255(p6842,p6844,p7052,p7053);
FA fa2271(p6846,p6848,p6862,p7054,p7055);
FA fa2272(p6864,p6868,p7023,p7056,p7057);
HA ha1256(p7025,p7027,p7058,p7059);
FA fa2273(p7035,p7041,p6852,p7060,p7061);
FA fa2274(p6854,p6856,p6878,p7062,p7063);
HA ha1257(p6880,p6884,p7064,p7065);
FA fa2275(p7031,p7033,p7037,p7066,p7067);
FA fa2276(p7039,p7051,p7053,p7068,p7069);
FA fa2277(p7059,p6860,p6866,p7070,p7071);
FA fa2278(p6870,p6872,p6874,p7072,p7073);
HA ha1258(p7043,p7045,p7074,p7075);
FA fa2279(p7047,p7049,p7055,p7076,p7077);
FA fa2280(p7057,p7061,p7065,p7078,p7079);
FA fa2281(p6876,p6882,p6886,p7080,p7081);
FA fa2282(p6888,p6890,p6902,p7082,p7083);
HA ha1259(p6908,p6910,p7084,p7085);
HA ha1260(p7063,p7067,p7086,p7087);
HA ha1261(p7069,p7075,p7088,p7089);
FA fa2283(p6892,p6894,p6896,p7090,p7091);
HA ha1262(p6898,p6900,p7092,p7093);
HA ha1263(p7071,p7073,p7094,p7095);
FA fa2284(p7077,p7079,p7085,p7096,p7097);
FA fa2285(p7087,p7089,p6904,p7098,p7099);
FA fa2286(p6906,p7081,p7083,p7100,p7101);
FA fa2287(p7093,p7095,p6912,p7102,p7103);
FA fa2288(p6914,p6916,p6918,p7104,p7105);
FA fa2289(p6920,p6922,p6928,p7106,p7107);
HA ha1264(p6930,p7091,p7108,p7109);
FA fa2290(p7097,p7099,p6924,p7110,p7111);
FA fa2291(p6926,p6938,p7101,p7112,p7113);
FA fa2292(p7103,p7109,p6932,p7114,p7115);
HA ha1265(p6934,p7105,p7116,p7117);
FA fa2293(p7107,p7111,p6936,p7118,p7119);
FA fa2294(p6940,p6948,p7113,p7120,p7121);
FA fa2295(p7115,p7117,p6942,p7122,p7123);
FA fa2296(p6944,p6946,p7119,p7124,p7125);
HA ha1266(p6950,p6956,p7126,p7127);
FA fa2297(p6958,p7121,p7123,p7128,p7129);
HA ha1267(p6952,p6954,p7130,p7131);
FA fa2298(p7125,p7127,p7129,p7132,p7133);
FA fa2299(p7131,p6960,p6962,p7134,p7135);
HA ha1268(p6964,p7133,p7136,p7137);
FA fa2300(p7137,p7135,p6966,p7138,p7139);
HA ha1269(p6968,p6970,p7140,p7141);
FA fa2301(p7139,p7141,p6972,p7142,p7143);
HA ha1270(p7143,p6974,p7144,p7145);
FA fa2302(ip_8_63,ip_9_62,ip_10_61,p7146,p7147);
HA ha1271(ip_11_60,ip_12_59,p7148,p7149);
FA fa2303(ip_13_58,ip_14_57,ip_15_56,p7150,p7151);
HA ha1272(ip_16_55,ip_17_54,p7152,p7153);
FA fa2304(ip_18_53,ip_19_52,ip_20_51,p7154,p7155);
FA fa2305(ip_21_50,ip_22_49,ip_23_48,p7156,p7157);
HA ha1273(ip_24_47,ip_25_46,p7158,p7159);
HA ha1274(ip_26_45,ip_27_44,p7160,p7161);
FA fa2306(ip_28_43,ip_29_42,ip_30_41,p7162,p7163);
FA fa2307(ip_31_40,ip_32_39,ip_33_38,p7164,p7165);
FA fa2308(ip_34_37,ip_35_36,ip_36_35,p7166,p7167);
FA fa2309(ip_37_34,ip_38_33,ip_39_32,p7168,p7169);
HA ha1275(ip_40_31,ip_41_30,p7170,p7171);
HA ha1276(ip_42_29,ip_43_28,p7172,p7173);
FA fa2310(ip_44_27,ip_45_26,ip_46_25,p7174,p7175);
FA fa2311(ip_47_24,ip_48_23,ip_49_22,p7176,p7177);
FA fa2312(ip_50_21,ip_51_20,ip_52_19,p7178,p7179);
FA fa2313(ip_53_18,ip_54_17,ip_55_16,p7180,p7181);
FA fa2314(ip_56_15,ip_57_14,ip_58_13,p7182,p7183);
FA fa2315(ip_59_12,ip_60_11,ip_61_10,p7184,p7185);
FA fa2316(ip_62_9,ip_63_8,p6978,p7186,p7187);
FA fa2317(p6984,p6988,p6994,p7188,p7189);
HA ha1277(p6998,p7000,p7190,p7191);
HA ha1278(p7012,p7014,p7192,p7193);
FA fa2318(p7149,p7153,p7159,p7194,p7195);
FA fa2319(p7161,p7171,p7173,p7196,p7197);
FA fa2320(p7028,p7147,p7151,p7198,p7199);
FA fa2321(p7155,p7157,p7163,p7200,p7201);
HA ha1279(p7165,p7167,p7202,p7203);
HA ha1280(p7169,p7175,p7204,p7205);
FA fa2322(p7177,p7179,p7181,p7206,p7207);
HA ha1281(p7183,p7185,p7208,p7209);
FA fa2323(p7187,p7191,p7193,p7210,p7211);
FA fa2324(p6980,p6982,p6986,p7212,p7213);
FA fa2325(p6990,p6992,p6996,p7214,p7215);
HA ha1282(p7002,p7004,p7216,p7217);
FA fa2326(p7006,p7008,p7010,p7218,p7219);
HA ha1283(p7016,p7018,p7220,p7221);
HA ha1284(p7020,p7034,p7222,p7223);
HA ha1285(p7040,p7189,p7224,p7225);
FA fa2327(p7195,p7197,p7203,p7226,p7227);
HA ha1286(p7205,p7209,p7228,p7229);
FA fa2328(p7022,p7024,p7026,p7230,p7231);
FA fa2329(p7050,p7052,p7058,p7232,p7233);
FA fa2330(p7199,p7201,p7207,p7234,p7235);
HA ha1287(p7211,p7217,p7236,p7237);
FA fa2331(p7221,p7223,p7225,p7238,p7239);
HA ha1288(p7229,p7030,p7240,p7241);
FA fa2332(p7032,p7036,p7038,p7242,p7243);
FA fa2333(p7064,p7213,p7215,p7244,p7245);
FA fa2334(p7219,p7227,p7237,p7246,p7247);
FA fa2335(p7042,p7044,p7046,p7248,p7249);
HA ha1289(p7048,p7054,p7250,p7251);
FA fa2336(p7056,p7060,p7074,p7252,p7253);
HA ha1290(p7231,p7233,p7254,p7255);
FA fa2337(p7235,p7239,p7241,p7256,p7257);
FA fa2338(p7062,p7066,p7068,p7258,p7259);
FA fa2339(p7084,p7086,p7088,p7260,p7261);
FA fa2340(p7243,p7245,p7247,p7262,p7263);
HA ha1291(p7251,p7255,p7264,p7265);
HA ha1292(p7070,p7072,p7266,p7267);
HA ha1293(p7076,p7078,p7268,p7269);
FA fa2341(p7092,p7094,p7249,p7270,p7271);
HA ha1294(p7253,p7257,p7272,p7273);
FA fa2342(p7265,p7080,p7082,p7274,p7275);
FA fa2343(p7259,p7261,p7263,p7276,p7277);
FA fa2344(p7267,p7269,p7273,p7278,p7279);
HA ha1295(p7090,p7096,p7280,p7281);
FA fa2345(p7098,p7108,p7271,p7282,p7283);
HA ha1296(p7100,p7102,p7284,p7285);
HA ha1297(p7275,p7277,p7286,p7287);
FA fa2346(p7279,p7281,p7104,p7288,p7289);
HA ha1298(p7106,p7110,p7290,p7291);
FA fa2347(p7116,p7283,p7285,p7292,p7293);
FA fa2348(p7287,p7112,p7114,p7294,p7295);
FA fa2349(p7289,p7291,p7118,p7296,p7297);
HA ha1299(p7293,p7120,p7298,p7299);
FA fa2350(p7122,p7126,p7295,p7300,p7301);
HA ha1300(p7297,p7124,p7302,p7303);
HA ha1301(p7130,p7299,p7304,p7305);
HA ha1302(p7128,p7301,p7306,p7307);
FA fa2351(p7303,p7305,p7132,p7308,p7309);
HA ha1303(p7136,p7307,p7310,p7311);
FA fa2352(p7309,p7311,p7134,p7312,p7313);
HA ha1304(p7313,p7138,p7314,p7315);
HA ha1305(p7140,p7315,p7316,p7317);
FA fa2353(p7317,p7142,p7144,p7318,p7319);
FA fa2354(ip_9_63,ip_10_62,ip_11_61,p7320,p7321);
HA ha1306(ip_12_60,ip_13_59,p7322,p7323);
HA ha1307(ip_14_58,ip_15_57,p7324,p7325);
HA ha1308(ip_16_56,ip_17_55,p7326,p7327);
HA ha1309(ip_18_54,ip_19_53,p7328,p7329);
FA fa2355(ip_20_52,ip_21_51,ip_22_50,p7330,p7331);
HA ha1310(ip_23_49,ip_24_48,p7332,p7333);
FA fa2356(ip_25_47,ip_26_46,ip_27_45,p7334,p7335);
HA ha1311(ip_28_44,ip_29_43,p7336,p7337);
HA ha1312(ip_30_42,ip_31_41,p7338,p7339);
HA ha1313(ip_32_40,ip_33_39,p7340,p7341);
HA ha1314(ip_34_38,ip_35_37,p7342,p7343);
FA fa2357(ip_36_36,ip_37_35,ip_38_34,p7344,p7345);
FA fa2358(ip_39_33,ip_40_32,ip_41_31,p7346,p7347);
FA fa2359(ip_42_30,ip_43_29,ip_44_28,p7348,p7349);
FA fa2360(ip_45_27,ip_46_26,ip_47_25,p7350,p7351);
FA fa2361(ip_48_24,ip_49_23,ip_50_22,p7352,p7353);
FA fa2362(ip_51_21,ip_52_20,ip_53_19,p7354,p7355);
FA fa2363(ip_54_18,ip_55_17,ip_56_16,p7356,p7357);
FA fa2364(ip_57_15,ip_58_14,ip_59_13,p7358,p7359);
FA fa2365(ip_60_12,ip_61_11,ip_62_10,p7360,p7361);
FA fa2366(ip_63_9,p7148,p7152,p7362,p7363);
FA fa2367(p7158,p7160,p7170,p7364,p7365);
FA fa2368(p7172,p7323,p7325,p7366,p7367);
HA ha1315(p7327,p7329,p7368,p7369);
HA ha1316(p7333,p7337,p7370,p7371);
HA ha1317(p7339,p7341,p7372,p7373);
FA fa2369(p7343,p7190,p7192,p7374,p7375);
HA ha1318(p7321,p7331,p7376,p7377);
FA fa2370(p7335,p7345,p7347,p7378,p7379);
FA fa2371(p7349,p7351,p7353,p7380,p7381);
FA fa2372(p7355,p7357,p7359,p7382,p7383);
HA ha1319(p7361,p7369,p7384,p7385);
HA ha1320(p7371,p7373,p7386,p7387);
FA fa2373(p7146,p7150,p7154,p7388,p7389);
HA ha1321(p7156,p7162,p7390,p7391);
FA fa2374(p7164,p7166,p7168,p7392,p7393);
HA ha1322(p7174,p7176,p7394,p7395);
HA ha1323(p7178,p7180,p7396,p7397);
FA fa2375(p7182,p7184,p7186,p7398,p7399);
FA fa2376(p7202,p7204,p7208,p7400,p7401);
FA fa2377(p7363,p7365,p7367,p7402,p7403);
HA ha1324(p7377,p7385,p7404,p7405);
FA fa2378(p7387,p7188,p7194,p7406,p7407);
FA fa2379(p7196,p7216,p7220,p7408,p7409);
FA fa2380(p7222,p7224,p7228,p7410,p7411);
HA ha1325(p7375,p7379,p7412,p7413);
FA fa2381(p7381,p7383,p7391,p7414,p7415);
HA ha1326(p7395,p7397,p7416,p7417);
FA fa2382(p7405,p7198,p7200,p7418,p7419);
HA ha1327(p7206,p7210,p7420,p7421);
FA fa2383(p7236,p7389,p7393,p7422,p7423);
FA fa2384(p7399,p7401,p7403,p7424,p7425);
FA fa2385(p7413,p7417,p7212,p7426,p7427);
FA fa2386(p7214,p7218,p7226,p7428,p7429);
FA fa2387(p7240,p7407,p7409,p7430,p7431);
FA fa2388(p7411,p7415,p7421,p7432,p7433);
FA fa2389(p7230,p7232,p7234,p7434,p7435);
FA fa2390(p7238,p7250,p7254,p7436,p7437);
FA fa2391(p7419,p7423,p7425,p7438,p7439);
FA fa2392(p7427,p7242,p7244,p7440,p7441);
FA fa2393(p7246,p7264,p7429,p7442,p7443);
HA ha1328(p7431,p7433,p7444,p7445);
FA fa2394(p7248,p7252,p7256,p7446,p7447);
FA fa2395(p7266,p7268,p7272,p7448,p7449);
FA fa2396(p7435,p7437,p7439,p7450,p7451);
HA ha1329(p7445,p7258,p7452,p7453);
FA fa2397(p7260,p7262,p7441,p7454,p7455);
HA ha1330(p7443,p7270,p7456,p7457);
FA fa2398(p7280,p7447,p7449,p7458,p7459);
HA ha1331(p7451,p7453,p7460,p7461);
HA ha1332(p7274,p7276,p7462,p7463);
FA fa2399(p7278,p7284,p7286,p7464,p7465);
HA ha1333(p7455,p7457,p7466,p7467);
FA fa2400(p7461,p7282,p7290,p7468,p7469);
FA fa2401(p7459,p7463,p7467,p7470,p7471);
HA ha1334(p7288,p7465,p7472,p7473);
FA fa2402(p7292,p7469,p7471,p7474,p7475);
FA fa2403(p7473,p7294,p7296,p7476,p7477);
FA fa2404(p7298,p7302,p7304,p7478,p7479);
HA ha1335(p7475,p7300,p7480,p7481);
HA ha1336(p7306,p7477,p7482,p7483);
HA ha1337(p7310,p7479,p7484,p7485);
FA fa2405(p7481,p7483,p7308,p7486,p7487);
FA fa2406(p7485,p7487,p7312,p7488,p7489);
FA fa2407(p7314,p7489,p7316,p7490,p7491);
HA ha1338(ip_10_63,ip_11_62,p7492,p7493);
FA fa2408(ip_12_61,ip_13_60,ip_14_59,p7494,p7495);
FA fa2409(ip_15_58,ip_16_57,ip_17_56,p7496,p7497);
HA ha1339(ip_18_55,ip_19_54,p7498,p7499);
FA fa2410(ip_20_53,ip_21_52,ip_22_51,p7500,p7501);
FA fa2411(ip_23_50,ip_24_49,ip_25_48,p7502,p7503);
FA fa2412(ip_26_47,ip_27_46,ip_28_45,p7504,p7505);
FA fa2413(ip_29_44,ip_30_43,ip_31_42,p7506,p7507);
HA ha1340(ip_32_41,ip_33_40,p7508,p7509);
FA fa2414(ip_34_39,ip_35_38,ip_36_37,p7510,p7511);
HA ha1341(ip_37_36,ip_38_35,p7512,p7513);
FA fa2415(ip_39_34,ip_40_33,ip_41_32,p7514,p7515);
FA fa2416(ip_42_31,ip_43_30,ip_44_29,p7516,p7517);
FA fa2417(ip_45_28,ip_46_27,ip_47_26,p7518,p7519);
FA fa2418(ip_48_25,ip_49_24,ip_50_23,p7520,p7521);
HA ha1342(ip_51_22,ip_52_21,p7522,p7523);
FA fa2419(ip_53_20,ip_54_19,ip_55_18,p7524,p7525);
FA fa2420(ip_56_17,ip_57_16,ip_58_15,p7526,p7527);
FA fa2421(ip_59_14,ip_60_13,ip_61_12,p7528,p7529);
HA ha1343(ip_62_11,ip_63_10,p7530,p7531);
HA ha1344(p7322,p7324,p7532,p7533);
HA ha1345(p7326,p7328,p7534,p7535);
FA fa2422(p7332,p7336,p7338,p7536,p7537);
FA fa2423(p7340,p7342,p7493,p7538,p7539);
FA fa2424(p7499,p7509,p7513,p7540,p7541);
FA fa2425(p7523,p7531,p7368,p7542,p7543);
FA fa2426(p7370,p7372,p7495,p7544,p7545);
HA ha1346(p7497,p7501,p7546,p7547);
FA fa2427(p7503,p7505,p7507,p7548,p7549);
HA ha1347(p7511,p7515,p7550,p7551);
FA fa2428(p7517,p7519,p7521,p7552,p7553);
FA fa2429(p7525,p7527,p7529,p7554,p7555);
FA fa2430(p7533,p7535,p7320,p7556,p7557);
FA fa2431(p7330,p7334,p7344,p7558,p7559);
HA ha1348(p7346,p7348,p7560,p7561);
HA ha1349(p7350,p7352,p7562,p7563);
FA fa2432(p7354,p7356,p7358,p7564,p7565);
FA fa2433(p7360,p7376,p7384,p7566,p7567);
HA ha1350(p7386,p7537,p7568,p7569);
HA ha1351(p7539,p7541,p7570,p7571);
HA ha1352(p7543,p7547,p7572,p7573);
HA ha1353(p7551,p7362,p7574,p7575);
FA fa2434(p7364,p7366,p7390,p7576,p7577);
FA fa2435(p7394,p7396,p7404,p7578,p7579);
HA ha1354(p7545,p7549,p7580,p7581);
FA fa2436(p7553,p7555,p7557,p7582,p7583);
HA ha1355(p7561,p7563,p7584,p7585);
HA ha1356(p7569,p7571,p7586,p7587);
HA ha1357(p7573,p7374,p7588,p7589);
FA fa2437(p7378,p7380,p7382,p7590,p7591);
FA fa2438(p7412,p7416,p7559,p7592,p7593);
HA ha1358(p7565,p7567,p7594,p7595);
FA fa2439(p7575,p7581,p7585,p7596,p7597);
FA fa2440(p7587,p7388,p7392,p7598,p7599);
HA ha1359(p7398,p7400,p7600,p7601);
HA ha1360(p7402,p7420,p7602,p7603);
HA ha1361(p7577,p7579,p7604,p7605);
FA fa2441(p7583,p7589,p7595,p7606,p7607);
FA fa2442(p7406,p7408,p7410,p7608,p7609);
HA ha1362(p7414,p7591,p7610,p7611);
FA fa2443(p7593,p7597,p7601,p7612,p7613);
FA fa2444(p7603,p7605,p7418,p7614,p7615);
FA fa2445(p7422,p7424,p7426,p7616,p7617);
FA fa2446(p7599,p7607,p7611,p7618,p7619);
FA fa2447(p7428,p7430,p7432,p7620,p7621);
FA fa2448(p7444,p7609,p7613,p7622,p7623);
HA ha1363(p7615,p7434,p7624,p7625);
HA ha1364(p7436,p7438,p7626,p7627);
FA fa2449(p7617,p7619,p7440,p7628,p7629);
FA fa2450(p7442,p7452,p7621,p7630,p7631);
FA fa2451(p7623,p7625,p7627,p7632,p7633);
FA fa2452(p7446,p7448,p7450,p7634,p7635);
FA fa2453(p7456,p7460,p7629,p7636,p7637);
HA ha1365(p7454,p7462,p7638,p7639);
HA ha1366(p7466,p7631,p7640,p7641);
FA fa2454(p7633,p7458,p7635,p7642,p7643);
HA ha1367(p7637,p7639,p7644,p7645);
HA ha1368(p7641,p7464,p7646,p7647);
HA ha1369(p7472,p7645,p7648,p7649);
HA ha1370(p7468,p7470,p7650,p7651);
FA fa2455(p7643,p7647,p7649,p7652,p7653);
HA ha1371(p7651,p7474,p7654,p7655);
FA fa2456(p7653,p7476,p7480,p7656,p7657);
HA ha1372(p7482,p7655,p7658,p7659);
FA fa2457(p7478,p7484,p7659,p7660,p7661);
FA fa2458(p7657,p7486,p7661,p7662,p7663);
FA fa2459(p7488,p7663,p7490,p7664,p7665);
HA ha1373(ip_11_63,ip_12_62,p7666,p7667);
FA fa2460(ip_13_61,ip_14_60,ip_15_59,p7668,p7669);
HA ha1374(ip_16_58,ip_17_57,p7670,p7671);
FA fa2461(ip_18_56,ip_19_55,ip_20_54,p7672,p7673);
FA fa2462(ip_21_53,ip_22_52,ip_23_51,p7674,p7675);
FA fa2463(ip_24_50,ip_25_49,ip_26_48,p7676,p7677);
HA ha1375(ip_27_47,ip_28_46,p7678,p7679);
FA fa2464(ip_29_45,ip_30_44,ip_31_43,p7680,p7681);
FA fa2465(ip_32_42,ip_33_41,ip_34_40,p7682,p7683);
HA ha1376(ip_35_39,ip_36_38,p7684,p7685);
HA ha1377(ip_37_37,ip_38_36,p7686,p7687);
FA fa2466(ip_39_35,ip_40_34,ip_41_33,p7688,p7689);
FA fa2467(ip_42_32,ip_43_31,ip_44_30,p7690,p7691);
FA fa2468(ip_45_29,ip_46_28,ip_47_27,p7692,p7693);
HA ha1378(ip_48_26,ip_49_25,p7694,p7695);
HA ha1379(ip_50_24,ip_51_23,p7696,p7697);
HA ha1380(ip_52_22,ip_53_21,p7698,p7699);
FA fa2469(ip_54_20,ip_55_19,ip_56_18,p7700,p7701);
HA ha1381(ip_57_17,ip_58_16,p7702,p7703);
FA fa2470(ip_59_15,ip_60_14,ip_61_13,p7704,p7705);
FA fa2471(ip_62_12,ip_63_11,p7492,p7706,p7707);
HA ha1382(p7498,p7508,p7708,p7709);
FA fa2472(p7512,p7522,p7530,p7710,p7711);
FA fa2473(p7667,p7671,p7679,p7712,p7713);
FA fa2474(p7685,p7687,p7695,p7714,p7715);
FA fa2475(p7697,p7699,p7703,p7716,p7717);
FA fa2476(p7532,p7534,p7669,p7718,p7719);
FA fa2477(p7673,p7675,p7677,p7720,p7721);
FA fa2478(p7681,p7683,p7689,p7722,p7723);
FA fa2479(p7691,p7693,p7701,p7724,p7725);
FA fa2480(p7705,p7707,p7709,p7726,p7727);
FA fa2481(p7494,p7496,p7500,p7728,p7729);
HA ha1383(p7502,p7504,p7730,p7731);
HA ha1384(p7506,p7510,p7732,p7733);
FA fa2482(p7514,p7516,p7518,p7734,p7735);
HA ha1385(p7520,p7524,p7736,p7737);
FA fa2483(p7526,p7528,p7546,p7738,p7739);
FA fa2484(p7550,p7711,p7713,p7740,p7741);
FA fa2485(p7715,p7717,p7536,p7742,p7743);
FA fa2486(p7538,p7540,p7542,p7744,p7745);
HA ha1386(p7560,p7562,p7746,p7747);
HA ha1387(p7568,p7570,p7748,p7749);
FA fa2487(p7572,p7719,p7721,p7750,p7751);
HA ha1388(p7723,p7725,p7752,p7753);
FA fa2488(p7727,p7731,p7733,p7754,p7755);
FA fa2489(p7737,p7544,p7548,p7756,p7757);
FA fa2490(p7552,p7554,p7556,p7758,p7759);
FA fa2491(p7574,p7580,p7584,p7760,p7761);
HA ha1389(p7586,p7729,p7762,p7763);
HA ha1390(p7735,p7739,p7764,p7765);
HA ha1391(p7741,p7743,p7766,p7767);
FA fa2492(p7747,p7749,p7753,p7768,p7769);
FA fa2493(p7558,p7564,p7566,p7770,p7771);
FA fa2494(p7588,p7594,p7745,p7772,p7773);
HA ha1392(p7751,p7755,p7774,p7775);
HA ha1393(p7763,p7765,p7776,p7777);
HA ha1394(p7767,p7576,p7778,p7779);
FA fa2495(p7578,p7582,p7600,p7780,p7781);
HA ha1395(p7602,p7604,p7782,p7783);
FA fa2496(p7757,p7759,p7761,p7784,p7785);
FA fa2497(p7769,p7775,p7777,p7786,p7787);
HA ha1396(p7590,p7592,p7788,p7789);
FA fa2498(p7596,p7610,p7771,p7790,p7791);
HA ha1397(p7773,p7779,p7792,p7793);
FA fa2499(p7783,p7598,p7606,p7794,p7795);
HA ha1398(p7781,p7785,p7796,p7797);
FA fa2500(p7787,p7789,p7793,p7798,p7799);
FA fa2501(p7608,p7612,p7614,p7800,p7801);
FA fa2502(p7791,p7797,p7616,p7802,p7803);
FA fa2503(p7618,p7624,p7626,p7804,p7805);
HA ha1399(p7795,p7799,p7806,p7807);
FA fa2504(p7620,p7622,p7801,p7808,p7809);
HA ha1400(p7803,p7807,p7810,p7811);
FA fa2505(p7628,p7805,p7811,p7812,p7813);
HA ha1401(p7630,p7632,p7814,p7815);
FA fa2506(p7638,p7640,p7809,p7816,p7817);
HA ha1402(p7634,p7636,p7818,p7819);
FA fa2507(p7644,p7813,p7815,p7820,p7821);
FA fa2508(p7646,p7648,p7817,p7822,p7823);
HA ha1403(p7819,p7642,p7824,p7825);
FA fa2509(p7650,p7821,p7823,p7826,p7827);
FA fa2510(p7825,p7652,p7654,p7828,p7829);
FA fa2511(p7827,p7658,p7829,p7830,p7831);
FA fa2512(p7656,p7831,p7660,p7832,p7833);
FA fa2513(p7833,p7662,p7664,p7834,p7835);
FA fa2514(ip_12_63,ip_13_62,ip_14_61,p7836,p7837);
FA fa2515(ip_15_60,ip_16_59,ip_17_58,p7838,p7839);
HA ha1404(ip_18_57,ip_19_56,p7840,p7841);
HA ha1405(ip_20_55,ip_21_54,p7842,p7843);
FA fa2516(ip_22_53,ip_23_52,ip_24_51,p7844,p7845);
FA fa2517(ip_25_50,ip_26_49,ip_27_48,p7846,p7847);
FA fa2518(ip_28_47,ip_29_46,ip_30_45,p7848,p7849);
FA fa2519(ip_31_44,ip_32_43,ip_33_42,p7850,p7851);
FA fa2520(ip_34_41,ip_35_40,ip_36_39,p7852,p7853);
FA fa2521(ip_37_38,ip_38_37,ip_39_36,p7854,p7855);
HA ha1406(ip_40_35,ip_41_34,p7856,p7857);
FA fa2522(ip_42_33,ip_43_32,ip_44_31,p7858,p7859);
FA fa2523(ip_45_30,ip_46_29,ip_47_28,p7860,p7861);
FA fa2524(ip_48_27,ip_49_26,ip_50_25,p7862,p7863);
HA ha1407(ip_51_24,ip_52_23,p7864,p7865);
FA fa2525(ip_53_22,ip_54_21,ip_55_20,p7866,p7867);
HA ha1408(ip_56_19,ip_57_18,p7868,p7869);
FA fa2526(ip_58_17,ip_59_16,ip_60_15,p7870,p7871);
FA fa2527(ip_61_14,ip_62_13,ip_63_12,p7872,p7873);
FA fa2528(p7666,p7670,p7678,p7874,p7875);
FA fa2529(p7684,p7686,p7694,p7876,p7877);
HA ha1409(p7696,p7698,p7878,p7879);
FA fa2530(p7702,p7841,p7843,p7880,p7881);
FA fa2531(p7857,p7865,p7869,p7882,p7883);
FA fa2532(p7708,p7837,p7839,p7884,p7885);
FA fa2533(p7845,p7847,p7849,p7886,p7887);
FA fa2534(p7851,p7853,p7855,p7888,p7889);
FA fa2535(p7859,p7861,p7863,p7890,p7891);
FA fa2536(p7867,p7871,p7873,p7892,p7893);
FA fa2537(p7879,p7668,p7672,p7894,p7895);
FA fa2538(p7674,p7676,p7680,p7896,p7897);
FA fa2539(p7682,p7688,p7690,p7898,p7899);
FA fa2540(p7692,p7700,p7704,p7900,p7901);
FA fa2541(p7706,p7875,p7877,p7902,p7903);
FA fa2542(p7881,p7883,p7710,p7904,p7905);
HA ha1410(p7712,p7714,p7906,p7907);
FA fa2543(p7716,p7730,p7732,p7908,p7909);
FA fa2544(p7736,p7885,p7887,p7910,p7911);
FA fa2545(p7889,p7891,p7893,p7912,p7913);
HA ha1411(p7718,p7720,p7914,p7915);
FA fa2546(p7722,p7724,p7726,p7916,p7917);
HA ha1412(p7746,p7748,p7918,p7919);
FA fa2547(p7752,p7895,p7897,p7920,p7921);
HA ha1413(p7899,p7901,p7922,p7923);
FA fa2548(p7903,p7905,p7907,p7924,p7925);
HA ha1414(p7728,p7734,p7926,p7927);
FA fa2549(p7738,p7740,p7742,p7928,p7929);
FA fa2550(p7762,p7764,p7766,p7930,p7931);
FA fa2551(p7909,p7911,p7913,p7932,p7933);
FA fa2552(p7915,p7919,p7923,p7934,p7935);
HA ha1415(p7744,p7750,p7936,p7937);
HA ha1416(p7754,p7774,p7938,p7939);
HA ha1417(p7776,p7917,p7940,p7941);
FA fa2553(p7921,p7925,p7927,p7942,p7943);
HA ha1418(p7756,p7758,p7944,p7945);
HA ha1419(p7760,p7768,p7946,p7947);
FA fa2554(p7778,p7782,p7929,p7948,p7949);
FA fa2555(p7931,p7933,p7935,p7950,p7951);
FA fa2556(p7937,p7939,p7941,p7952,p7953);
FA fa2557(p7770,p7772,p7788,p7954,p7955);
FA fa2558(p7792,p7943,p7945,p7956,p7957);
FA fa2559(p7947,p7780,p7784,p7958,p7959);
HA ha1420(p7786,p7796,p7960,p7961);
FA fa2560(p7949,p7951,p7953,p7962,p7963);
FA fa2561(p7790,p7955,p7957,p7964,p7965);
HA ha1421(p7961,p7794,p7966,p7967);
FA fa2562(p7798,p7806,p7959,p7968,p7969);
HA ha1422(p7963,p7800,p7970,p7971);
FA fa2563(p7802,p7810,p7965,p7972,p7973);
FA fa2564(p7967,p7804,p7969,p7974,p7975);
FA fa2565(p7971,p7808,p7814,p7976,p7977);
HA ha1423(p7973,p7812,p7978,p7979);
FA fa2566(p7818,p7975,p7816,p7980,p7981);
FA fa2567(p7977,p7979,p7820,p7982,p7983);
FA fa2568(p7824,p7981,p7822,p7984,p7985);
FA fa2569(p7983,p7826,p7985,p7986,p7987);
FA fa2570(p7828,p7987,p7830,p7988,p7989);
HA ha1424(p7989,p7832,p7990,p7991);
HA ha1425(ip_13_63,ip_14_62,p7992,p7993);
HA ha1426(ip_15_61,ip_16_60,p7994,p7995);
FA fa2571(ip_17_59,ip_18_58,ip_19_57,p7996,p7997);
FA fa2572(ip_20_56,ip_21_55,ip_22_54,p7998,p7999);
HA ha1427(ip_23_53,ip_24_52,p8000,p8001);
FA fa2573(ip_25_51,ip_26_50,ip_27_49,p8002,p8003);
FA fa2574(ip_28_48,ip_29_47,ip_30_46,p8004,p8005);
FA fa2575(ip_31_45,ip_32_44,ip_33_43,p8006,p8007);
FA fa2576(ip_34_42,ip_35_41,ip_36_40,p8008,p8009);
HA ha1428(ip_37_39,ip_38_38,p8010,p8011);
HA ha1429(ip_39_37,ip_40_36,p8012,p8013);
FA fa2577(ip_41_35,ip_42_34,ip_43_33,p8014,p8015);
FA fa2578(ip_44_32,ip_45_31,ip_46_30,p8016,p8017);
HA ha1430(ip_47_29,ip_48_28,p8018,p8019);
HA ha1431(ip_49_27,ip_50_26,p8020,p8021);
FA fa2579(ip_51_25,ip_52_24,ip_53_23,p8022,p8023);
FA fa2580(ip_54_22,ip_55_21,ip_56_20,p8024,p8025);
FA fa2581(ip_57_19,ip_58_18,ip_59_17,p8026,p8027);
HA ha1432(ip_60_16,ip_61_15,p8028,p8029);
HA ha1433(ip_62_14,ip_63_13,p8030,p8031);
FA fa2582(p7840,p7842,p7856,p8032,p8033);
FA fa2583(p7864,p7868,p7993,p8034,p8035);
FA fa2584(p7995,p8001,p8011,p8036,p8037);
FA fa2585(p8013,p8019,p8021,p8038,p8039);
FA fa2586(p8029,p8031,p7878,p8040,p8041);
FA fa2587(p7997,p7999,p8003,p8042,p8043);
HA ha1434(p8005,p8007,p8044,p8045);
HA ha1435(p8009,p8015,p8046,p8047);
HA ha1436(p8017,p8023,p8048,p8049);
FA fa2588(p8025,p8027,p7836,p8050,p8051);
HA ha1437(p7838,p7844,p8052,p8053);
FA fa2589(p7846,p7848,p7850,p8054,p8055);
FA fa2590(p7852,p7854,p7858,p8056,p8057);
FA fa2591(p7860,p7862,p7866,p8058,p8059);
HA ha1438(p7870,p7872,p8060,p8061);
FA fa2592(p8033,p8035,p8037,p8062,p8063);
FA fa2593(p8039,p8041,p8045,p8064,p8065);
FA fa2594(p8047,p8049,p7874,p8066,p8067);
FA fa2595(p7876,p7880,p7882,p8068,p8069);
HA ha1439(p8043,p8051,p8070,p8071);
HA ha1440(p8053,p8061,p8072,p8073);
FA fa2596(p7884,p7886,p7888,p8074,p8075);
FA fa2597(p7890,p7892,p7906,p8076,p8077);
FA fa2598(p8055,p8057,p8059,p8078,p8079);
HA ha1441(p8063,p8065,p8080,p8081);
HA ha1442(p8067,p8071,p8082,p8083);
HA ha1443(p8073,p7894,p8084,p8085);
HA ha1444(p7896,p7898,p8086,p8087);
FA fa2599(p7900,p7902,p7904,p8088,p8089);
FA fa2600(p7914,p7918,p7922,p8090,p8091);
HA ha1445(p8069,p8081,p8092,p8093);
FA fa2601(p8083,p7908,p7910,p8094,p8095);
FA fa2602(p7912,p7926,p8075,p8096,p8097);
FA fa2603(p8077,p8079,p8085,p8098,p8099);
HA ha1446(p8087,p8093,p8100,p8101);
HA ha1447(p7916,p7920,p8102,p8103);
FA fa2604(p7924,p7936,p7938,p8104,p8105);
FA fa2605(p7940,p8089,p8091,p8106,p8107);
FA fa2606(p8101,p7928,p7930,p8108,p8109);
FA fa2607(p7932,p7934,p7944,p8110,p8111);
HA ha1448(p7946,p8095,p8112,p8113);
HA ha1449(p8097,p8099,p8114,p8115);
FA fa2608(p8103,p7942,p8105,p8116,p8117);
FA fa2609(p8107,p8113,p8115,p8118,p8119);
FA fa2610(p7948,p7950,p7952,p8120,p8121);
FA fa2611(p7960,p8109,p8111,p8122,p8123);
FA fa2612(p7954,p7956,p8117,p8124,p8125);
FA fa2613(p8119,p7958,p7962,p8126,p8127);
FA fa2614(p7966,p8121,p8123,p8128,p8129);
FA fa2615(p7964,p7970,p8125,p8130,p8131);
HA ha1450(p7968,p8127,p8132,p8133);
FA fa2616(p8129,p7972,p8131,p8134,p8135);
HA ha1451(p8133,p7974,p8136,p8137);
HA ha1452(p7978,p7976,p8138,p8139);
HA ha1453(p8135,p8137,p8140,p8141);
FA fa2617(p7980,p8139,p8141,p8142,p8143);
FA fa2618(p7982,p7984,p8143,p8144,p8145);
HA ha1454(p7986,p8145,p8146,p8147);
FA fa2619(p8147,p7988,p7990,p8148,p8149);
FA fa2620(ip_14_63,ip_15_62,ip_16_61,p8150,p8151);
FA fa2621(ip_17_60,ip_18_59,ip_19_58,p8152,p8153);
FA fa2622(ip_20_57,ip_21_56,ip_22_55,p8154,p8155);
FA fa2623(ip_23_54,ip_24_53,ip_25_52,p8156,p8157);
FA fa2624(ip_26_51,ip_27_50,ip_28_49,p8158,p8159);
HA ha1455(ip_29_48,ip_30_47,p8160,p8161);
HA ha1456(ip_31_46,ip_32_45,p8162,p8163);
FA fa2625(ip_33_44,ip_34_43,ip_35_42,p8164,p8165);
FA fa2626(ip_36_41,ip_37_40,ip_38_39,p8166,p8167);
FA fa2627(ip_39_38,ip_40_37,ip_41_36,p8168,p8169);
FA fa2628(ip_42_35,ip_43_34,ip_44_33,p8170,p8171);
HA ha1457(ip_45_32,ip_46_31,p8172,p8173);
FA fa2629(ip_47_30,ip_48_29,ip_49_28,p8174,p8175);
HA ha1458(ip_50_27,ip_51_26,p8176,p8177);
FA fa2630(ip_52_25,ip_53_24,ip_54_23,p8178,p8179);
HA ha1459(ip_55_22,ip_56_21,p8180,p8181);
FA fa2631(ip_57_20,ip_58_19,ip_59_18,p8182,p8183);
FA fa2632(ip_60_17,ip_61_16,ip_62_15,p8184,p8185);
FA fa2633(ip_63_14,p7992,p7994,p8186,p8187);
FA fa2634(p8000,p8010,p8012,p8188,p8189);
FA fa2635(p8018,p8020,p8028,p8190,p8191);
HA ha1460(p8030,p8161,p8192,p8193);
HA ha1461(p8163,p8173,p8194,p8195);
FA fa2636(p8177,p8181,p8151,p8196,p8197);
HA ha1462(p8153,p8155,p8198,p8199);
HA ha1463(p8157,p8159,p8200,p8201);
FA fa2637(p8165,p8167,p8169,p8202,p8203);
HA ha1464(p8171,p8175,p8204,p8205);
FA fa2638(p8179,p8183,p8185,p8206,p8207);
FA fa2639(p8193,p8195,p7996,p8208,p8209);
FA fa2640(p7998,p8002,p8004,p8210,p8211);
FA fa2641(p8006,p8008,p8014,p8212,p8213);
FA fa2642(p8016,p8022,p8024,p8214,p8215);
HA ha1465(p8026,p8044,p8216,p8217);
HA ha1466(p8046,p8048,p8218,p8219);
FA fa2643(p8187,p8189,p8191,p8220,p8221);
FA fa2644(p8197,p8199,p8201,p8222,p8223);
HA ha1467(p8205,p8032,p8224,p8225);
FA fa2645(p8034,p8036,p8038,p8226,p8227);
FA fa2646(p8040,p8052,p8060,p8228,p8229);
FA fa2647(p8203,p8207,p8209,p8230,p8231);
FA fa2648(p8217,p8219,p8042,p8232,p8233);
HA ha1468(p8050,p8070,p8234,p8235);
HA ha1469(p8072,p8211,p8236,p8237);
FA fa2649(p8213,p8215,p8221,p8238,p8239);
FA fa2650(p8223,p8225,p8054,p8240,p8241);
FA fa2651(p8056,p8058,p8062,p8242,p8243);
FA fa2652(p8064,p8066,p8080,p8244,p8245);
HA ha1470(p8082,p8227,p8246,p8247);
HA ha1471(p8229,p8231,p8248,p8249);
FA fa2653(p8233,p8235,p8237,p8250,p8251);
FA fa2654(p8068,p8084,p8086,p8252,p8253);
FA fa2655(p8092,p8239,p8241,p8254,p8255);
HA ha1472(p8247,p8249,p8256,p8257);
FA fa2656(p8074,p8076,p8078,p8258,p8259);
HA ha1473(p8100,p8243,p8260,p8261);
HA ha1474(p8245,p8251,p8262,p8263);
FA fa2657(p8257,p8088,p8090,p8264,p8265);
FA fa2658(p8102,p8253,p8255,p8266,p8267);
FA fa2659(p8261,p8263,p8094,p8268,p8269);
FA fa2660(p8096,p8098,p8112,p8270,p8271);
HA ha1475(p8114,p8259,p8272,p8273);
FA fa2661(p8104,p8106,p8265,p8274,p8275);
FA fa2662(p8267,p8269,p8273,p8276,p8277);
FA fa2663(p8108,p8110,p8271,p8278,p8279);
HA ha1476(p8116,p8118,p8280,p8281);
FA fa2664(p8275,p8277,p8120,p8282,p8283);
HA ha1477(p8122,p8279,p8284,p8285);
FA fa2665(p8281,p8124,p8283,p8286,p8287);
FA fa2666(p8285,p8126,p8128,p8288,p8289);
FA fa2667(p8132,p8130,p8287,p8290,p8291);
FA fa2668(p8136,p8289,p8134,p8292,p8293);
HA ha1478(p8138,p8140,p8294,p8295);
FA fa2669(p8291,p8293,p8295,p8296,p8297);
HA ha1479(p8142,p8297,p8298,p8299);
HA ha1480(p8299,p8144,p8300,p8301);
FA fa2670(p8146,p8301,p8148,p8302,p8303);
HA ha1481(ip_15_63,ip_16_62,p8304,p8305);
HA ha1482(ip_17_61,ip_18_60,p8306,p8307);
FA fa2671(ip_19_59,ip_20_58,ip_21_57,p8308,p8309);
FA fa2672(ip_22_56,ip_23_55,ip_24_54,p8310,p8311);
HA ha1483(ip_25_53,ip_26_52,p8312,p8313);
HA ha1484(ip_27_51,ip_28_50,p8314,p8315);
FA fa2673(ip_29_49,ip_30_48,ip_31_47,p8316,p8317);
HA ha1485(ip_32_46,ip_33_45,p8318,p8319);
FA fa2674(ip_34_44,ip_35_43,ip_36_42,p8320,p8321);
FA fa2675(ip_37_41,ip_38_40,ip_39_39,p8322,p8323);
FA fa2676(ip_40_38,ip_41_37,ip_42_36,p8324,p8325);
FA fa2677(ip_43_35,ip_44_34,ip_45_33,p8326,p8327);
FA fa2678(ip_46_32,ip_47_31,ip_48_30,p8328,p8329);
FA fa2679(ip_49_29,ip_50_28,ip_51_27,p8330,p8331);
HA ha1486(ip_52_26,ip_53_25,p8332,p8333);
FA fa2680(ip_54_24,ip_55_23,ip_56_22,p8334,p8335);
HA ha1487(ip_57_21,ip_58_20,p8336,p8337);
HA ha1488(ip_59_19,ip_60_18,p8338,p8339);
FA fa2681(ip_61_17,ip_62_16,ip_63_15,p8340,p8341);
HA ha1489(p8160,p8162,p8342,p8343);
FA fa2682(p8172,p8176,p8180,p8344,p8345);
FA fa2683(p8305,p8307,p8313,p8346,p8347);
FA fa2684(p8315,p8319,p8333,p8348,p8349);
HA ha1490(p8337,p8339,p8350,p8351);
FA fa2685(p8192,p8194,p8309,p8352,p8353);
FA fa2686(p8311,p8317,p8321,p8354,p8355);
FA fa2687(p8323,p8325,p8327,p8356,p8357);
FA fa2688(p8329,p8331,p8335,p8358,p8359);
HA ha1491(p8341,p8343,p8360,p8361);
FA fa2689(p8351,p8150,p8152,p8362,p8363);
FA fa2690(p8154,p8156,p8158,p8364,p8365);
FA fa2691(p8164,p8166,p8168,p8366,p8367);
HA ha1492(p8170,p8174,p8368,p8369);
HA ha1493(p8178,p8182,p8370,p8371);
HA ha1494(p8184,p8198,p8372,p8373);
HA ha1495(p8200,p8204,p8374,p8375);
HA ha1496(p8345,p8347,p8376,p8377);
FA fa2692(p8349,p8361,p8186,p8378,p8379);
FA fa2693(p8188,p8190,p8196,p8380,p8381);
HA ha1497(p8216,p8218,p8382,p8383);
FA fa2694(p8353,p8355,p8357,p8384,p8385);
FA fa2695(p8359,p8369,p8371,p8386,p8387);
FA fa2696(p8373,p8375,p8377,p8388,p8389);
FA fa2697(p8202,p8206,p8208,p8390,p8391);
FA fa2698(p8224,p8363,p8365,p8392,p8393);
FA fa2699(p8367,p8379,p8383,p8394,p8395);
HA ha1498(p8210,p8212,p8396,p8397);
FA fa2700(p8214,p8220,p8222,p8398,p8399);
FA fa2701(p8234,p8236,p8381,p8400,p8401);
FA fa2702(p8385,p8387,p8389,p8402,p8403);
FA fa2703(p8226,p8228,p8230,p8404,p8405);
FA fa2704(p8232,p8246,p8248,p8406,p8407);
FA fa2705(p8391,p8393,p8395,p8408,p8409);
FA fa2706(p8397,p8238,p8240,p8410,p8411);
HA ha1499(p8256,p8399,p8412,p8413);
HA ha1500(p8401,p8403,p8414,p8415);
HA ha1501(p8242,p8244,p8416,p8417);
FA fa2707(p8250,p8260,p8262,p8418,p8419);
FA fa2708(p8405,p8407,p8409,p8420,p8421);
HA ha1502(p8413,p8415,p8422,p8423);
FA fa2709(p8252,p8254,p8411,p8424,p8425);
HA ha1503(p8417,p8423,p8426,p8427);
HA ha1504(p8258,p8272,p8428,p8429);
FA fa2710(p8419,p8421,p8427,p8430,p8431);
FA fa2711(p8264,p8266,p8268,p8432,p8433);
HA ha1505(p8425,p8429,p8434,p8435);
HA ha1506(p8270,p8431,p8436,p8437);
FA fa2712(p8435,p8274,p8276,p8438,p8439);
FA fa2713(p8280,p8433,p8437,p8440,p8441);
FA fa2714(p8278,p8284,p8282,p8442,p8443);
FA fa2715(p8439,p8441,p8443,p8444,p8445);
HA ha1507(p8286,p8445,p8446,p8447);
HA ha1508(p8288,p8447,p8448,p8449);
FA fa2716(p8290,p8294,p8449,p8450,p8451);
FA fa2717(p8292,p8451,p8296,p8452,p8453);
HA ha1509(p8298,p8453,p8454,p8455);
FA fa2718(p8300,p8455,p8302,p8456,p8457);
FA fa2719(ip_16_63,ip_17_62,ip_18_61,p8458,p8459);
HA ha1510(ip_19_60,ip_20_59,p8460,p8461);
HA ha1511(ip_21_58,ip_22_57,p8462,p8463);
FA fa2720(ip_23_56,ip_24_55,ip_25_54,p8464,p8465);
FA fa2721(ip_26_53,ip_27_52,ip_28_51,p8466,p8467);
HA ha1512(ip_29_50,ip_30_49,p8468,p8469);
HA ha1513(ip_31_48,ip_32_47,p8470,p8471);
FA fa2722(ip_33_46,ip_34_45,ip_35_44,p8472,p8473);
HA ha1514(ip_36_43,ip_37_42,p8474,p8475);
FA fa2723(ip_38_41,ip_39_40,ip_40_39,p8476,p8477);
FA fa2724(ip_41_38,ip_42_37,ip_43_36,p8478,p8479);
FA fa2725(ip_44_35,ip_45_34,ip_46_33,p8480,p8481);
FA fa2726(ip_47_32,ip_48_31,ip_49_30,p8482,p8483);
HA ha1515(ip_50_29,ip_51_28,p8484,p8485);
FA fa2727(ip_52_27,ip_53_26,ip_54_25,p8486,p8487);
FA fa2728(ip_55_24,ip_56_23,ip_57_22,p8488,p8489);
FA fa2729(ip_58_21,ip_59_20,ip_60_19,p8490,p8491);
FA fa2730(ip_61_18,ip_62_17,ip_63_16,p8492,p8493);
FA fa2731(p8304,p8306,p8312,p8494,p8495);
HA ha1516(p8314,p8318,p8496,p8497);
FA fa2732(p8332,p8336,p8338,p8498,p8499);
HA ha1517(p8461,p8463,p8500,p8501);
FA fa2733(p8469,p8471,p8475,p8502,p8503);
FA fa2734(p8485,p8342,p8350,p8504,p8505);
HA ha1518(p8459,p8465,p8506,p8507);
HA ha1519(p8467,p8473,p8508,p8509);
FA fa2735(p8477,p8479,p8481,p8510,p8511);
HA ha1520(p8483,p8487,p8512,p8513);
HA ha1521(p8489,p8491,p8514,p8515);
FA fa2736(p8493,p8497,p8501,p8516,p8517);
FA fa2737(p8308,p8310,p8316,p8518,p8519);
FA fa2738(p8320,p8322,p8324,p8520,p8521);
FA fa2739(p8326,p8328,p8330,p8522,p8523);
FA fa2740(p8334,p8340,p8360,p8524,p8525);
FA fa2741(p8495,p8499,p8503,p8526,p8527);
HA ha1522(p8507,p8509,p8528,p8529);
FA fa2742(p8513,p8515,p8344,p8530,p8531);
FA fa2743(p8346,p8348,p8368,p8532,p8533);
FA fa2744(p8370,p8372,p8374,p8534,p8535);
HA ha1523(p8376,p8505,p8536,p8537);
FA fa2745(p8511,p8517,p8529,p8538,p8539);
HA ha1524(p8352,p8354,p8540,p8541);
HA ha1525(p8356,p8358,p8542,p8543);
FA fa2746(p8382,p8519,p8521,p8544,p8545);
HA ha1526(p8523,p8525,p8546,p8547);
FA fa2747(p8527,p8531,p8537,p8548,p8549);
FA fa2748(p8362,p8364,p8366,p8550,p8551);
HA ha1527(p8378,p8533,p8552,p8553);
HA ha1528(p8535,p8539,p8554,p8555);
FA fa2749(p8541,p8543,p8547,p8556,p8557);
FA fa2750(p8380,p8384,p8386,p8558,p8559);
FA fa2751(p8388,p8396,p8545,p8560,p8561);
FA fa2752(p8549,p8553,p8555,p8562,p8563);
FA fa2753(p8390,p8392,p8394,p8564,p8565);
FA fa2754(p8551,p8557,p8398,p8566,p8567);
HA ha1529(p8400,p8402,p8568,p8569);
HA ha1530(p8412,p8414,p8570,p8571);
FA fa2755(p8559,p8561,p8563,p8572,p8573);
HA ha1531(p8404,p8406,p8574,p8575);
HA ha1532(p8408,p8416,p8576,p8577);
FA fa2756(p8422,p8565,p8567,p8578,p8579);
FA fa2757(p8569,p8571,p8410,p8580,p8581);
FA fa2758(p8426,p8573,p8575,p8582,p8583);
HA ha1533(p8577,p8418,p8584,p8585);
HA ha1534(p8420,p8428,p8586,p8587);
FA fa2759(p8579,p8581,p8424,p8588,p8589);
HA ha1535(p8434,p8583,p8590,p8591);
FA fa2760(p8585,p8587,p8430,p8592,p8593);
FA fa2761(p8436,p8589,p8591,p8594,p8595);
HA ha1536(p8432,p8593,p8596,p8597);
FA fa2762(p8595,p8597,p8438,p8598,p8599);
FA fa2763(p8440,p8442,p8599,p8600,p8601);
HA ha1537(p8444,p8446,p8602,p8603);
FA fa2764(p8448,p8601,p8603,p8604,p8605);
FA fa2765(p8605,p8450,p8452,p8606,p8607);
FA fa2766(p8454,p8607,p8456,p8608,p8609);
FA fa2767(ip_17_63,ip_18_62,ip_19_61,p8610,p8611);
HA ha1538(ip_20_60,ip_21_59,p8612,p8613);
FA fa2768(ip_22_58,ip_23_57,ip_24_56,p8614,p8615);
FA fa2769(ip_25_55,ip_26_54,ip_27_53,p8616,p8617);
FA fa2770(ip_28_52,ip_29_51,ip_30_50,p8618,p8619);
FA fa2771(ip_31_49,ip_32_48,ip_33_47,p8620,p8621);
HA ha1539(ip_34_46,ip_35_45,p8622,p8623);
HA ha1540(ip_36_44,ip_37_43,p8624,p8625);
FA fa2772(ip_38_42,ip_39_41,ip_40_40,p8626,p8627);
HA ha1541(ip_41_39,ip_42_38,p8628,p8629);
FA fa2773(ip_43_37,ip_44_36,ip_45_35,p8630,p8631);
FA fa2774(ip_46_34,ip_47_33,ip_48_32,p8632,p8633);
HA ha1542(ip_49_31,ip_50_30,p8634,p8635);
HA ha1543(ip_51_29,ip_52_28,p8636,p8637);
FA fa2775(ip_53_27,ip_54_26,ip_55_25,p8638,p8639);
FA fa2776(ip_56_24,ip_57_23,ip_58_22,p8640,p8641);
HA ha1544(ip_59_21,ip_60_20,p8642,p8643);
FA fa2777(ip_61_19,ip_62_18,ip_63_17,p8644,p8645);
HA ha1545(p8460,p8462,p8646,p8647);
FA fa2778(p8468,p8470,p8474,p8648,p8649);
FA fa2779(p8484,p8613,p8623,p8650,p8651);
HA ha1546(p8625,p8629,p8652,p8653);
HA ha1547(p8635,p8637,p8654,p8655);
HA ha1548(p8643,p8496,p8656,p8657);
FA fa2780(p8500,p8611,p8615,p8658,p8659);
FA fa2781(p8617,p8619,p8621,p8660,p8661);
HA ha1549(p8627,p8631,p8662,p8663);
HA ha1550(p8633,p8639,p8664,p8665);
FA fa2782(p8641,p8645,p8647,p8666,p8667);
HA ha1551(p8653,p8655,p8668,p8669);
HA ha1552(p8458,p8464,p8670,p8671);
FA fa2783(p8466,p8472,p8476,p8672,p8673);
HA ha1553(p8478,p8480,p8674,p8675);
FA fa2784(p8482,p8486,p8488,p8676,p8677);
FA fa2785(p8490,p8492,p8506,p8678,p8679);
HA ha1554(p8508,p8512,p8680,p8681);
FA fa2786(p8514,p8649,p8651,p8682,p8683);
FA fa2787(p8657,p8663,p8665,p8684,p8685);
FA fa2788(p8669,p8494,p8498,p8686,p8687);
HA ha1555(p8502,p8528,p8688,p8689);
HA ha1556(p8659,p8661,p8690,p8691);
FA fa2789(p8667,p8671,p8675,p8692,p8693);
HA ha1557(p8681,p8504,p8694,p8695);
HA ha1558(p8510,p8516,p8696,p8697);
HA ha1559(p8536,p8673,p8698,p8699);
HA ha1560(p8677,p8679,p8700,p8701);
FA fa2790(p8683,p8685,p8689,p8702,p8703);
FA fa2791(p8691,p8518,p8520,p8704,p8705);
FA fa2792(p8522,p8524,p8526,p8706,p8707);
FA fa2793(p8530,p8540,p8542,p8708,p8709);
FA fa2794(p8546,p8687,p8693,p8710,p8711);
FA fa2795(p8695,p8697,p8699,p8712,p8713);
HA ha1561(p8701,p8532,p8714,p8715);
HA ha1562(p8534,p8538,p8716,p8717);
FA fa2796(p8552,p8554,p8703,p8718,p8719);
FA fa2797(p8544,p8548,p8705,p8720,p8721);
FA fa2798(p8707,p8709,p8711,p8722,p8723);
FA fa2799(p8713,p8715,p8717,p8724,p8725);
FA fa2800(p8550,p8556,p8719,p8726,p8727);
FA fa2801(p8558,p8560,p8562,p8728,p8729);
FA fa2802(p8568,p8570,p8721,p8730,p8731);
HA ha1563(p8723,p8725,p8732,p8733);
HA ha1564(p8564,p8566,p8734,p8735);
FA fa2803(p8574,p8576,p8727,p8736,p8737);
FA fa2804(p8733,p8572,p8729,p8738,p8739);
HA ha1565(p8731,p8735,p8740,p8741);
FA fa2805(p8578,p8580,p8584,p8742,p8743);
FA fa2806(p8586,p8737,p8741,p8744,p8745);
FA fa2807(p8582,p8590,p8739,p8746,p8747);
FA fa2808(p8588,p8743,p8745,p8748,p8749);
HA ha1566(p8592,p8596,p8750,p8751);
FA fa2809(p8747,p8594,p8749,p8752,p8753);
FA fa2810(p8751,p8598,p8753,p8754,p8755);
FA fa2811(p8602,p8600,p8755,p8756,p8757);
FA fa2812(p8604,p8757,p8606,p8758,p8759);
FA fa2813(ip_18_63,ip_19_62,ip_20_61,p8760,p8761);
FA fa2814(ip_21_60,ip_22_59,ip_23_58,p8762,p8763);
FA fa2815(ip_24_57,ip_25_56,ip_26_55,p8764,p8765);
HA ha1567(ip_27_54,ip_28_53,p8766,p8767);
FA fa2816(ip_29_52,ip_30_51,ip_31_50,p8768,p8769);
FA fa2817(ip_32_49,ip_33_48,ip_34_47,p8770,p8771);
HA ha1568(ip_35_46,ip_36_45,p8772,p8773);
HA ha1569(ip_37_44,ip_38_43,p8774,p8775);
HA ha1570(ip_39_42,ip_40_41,p8776,p8777);
HA ha1571(ip_41_40,ip_42_39,p8778,p8779);
HA ha1572(ip_43_38,ip_44_37,p8780,p8781);
FA fa2818(ip_45_36,ip_46_35,ip_47_34,p8782,p8783);
FA fa2819(ip_48_33,ip_49_32,ip_50_31,p8784,p8785);
FA fa2820(ip_51_30,ip_52_29,ip_53_28,p8786,p8787);
HA ha1573(ip_54_27,ip_55_26,p8788,p8789);
HA ha1574(ip_56_25,ip_57_24,p8790,p8791);
FA fa2821(ip_58_23,ip_59_22,ip_60_21,p8792,p8793);
HA ha1575(ip_61_20,ip_62_19,p8794,p8795);
FA fa2822(ip_63_18,p8612,p8622,p8796,p8797);
FA fa2823(p8624,p8628,p8634,p8798,p8799);
FA fa2824(p8636,p8642,p8767,p8800,p8801);
HA ha1576(p8773,p8775,p8802,p8803);
HA ha1577(p8777,p8779,p8804,p8805);
FA fa2825(p8781,p8789,p8791,p8806,p8807);
FA fa2826(p8795,p8646,p8652,p8808,p8809);
FA fa2827(p8654,p8761,p8763,p8810,p8811);
FA fa2828(p8765,p8769,p8771,p8812,p8813);
HA ha1578(p8783,p8785,p8814,p8815);
FA fa2829(p8787,p8793,p8803,p8816,p8817);
FA fa2830(p8805,p8610,p8614,p8818,p8819);
FA fa2831(p8616,p8618,p8620,p8820,p8821);
FA fa2832(p8626,p8630,p8632,p8822,p8823);
FA fa2833(p8638,p8640,p8644,p8824,p8825);
FA fa2834(p8656,p8662,p8664,p8826,p8827);
FA fa2835(p8668,p8797,p8799,p8828,p8829);
FA fa2836(p8801,p8807,p8815,p8830,p8831);
FA fa2837(p8648,p8650,p8670,p8832,p8833);
HA ha1579(p8674,p8680,p8834,p8835);
HA ha1580(p8809,p8811,p8836,p8837);
FA fa2838(p8813,p8817,p8658,p8838,p8839);
FA fa2839(p8660,p8666,p8688,p8840,p8841);
FA fa2840(p8690,p8819,p8821,p8842,p8843);
HA ha1581(p8823,p8825,p8844,p8845);
HA ha1582(p8827,p8829,p8846,p8847);
FA fa2841(p8831,p8835,p8837,p8848,p8849);
HA ha1583(p8672,p8676,p8850,p8851);
FA fa2842(p8678,p8682,p8684,p8852,p8853);
FA fa2843(p8694,p8696,p8698,p8854,p8855);
FA fa2844(p8700,p8833,p8839,p8856,p8857);
FA fa2845(p8845,p8847,p8686,p8858,p8859);
FA fa2846(p8692,p8841,p8843,p8860,p8861);
HA ha1584(p8849,p8851,p8862,p8863);
FA fa2847(p8702,p8714,p8716,p8864,p8865);
FA fa2848(p8853,p8855,p8857,p8866,p8867);
FA fa2849(p8859,p8863,p8704,p8868,p8869);
FA fa2850(p8706,p8708,p8710,p8870,p8871);
HA ha1585(p8712,p8861,p8872,p8873);
FA fa2851(p8718,p8865,p8867,p8874,p8875);
HA ha1586(p8869,p8873,p8876,p8877);
HA ha1587(p8720,p8722,p8878,p8879);
FA fa2852(p8724,p8732,p8871,p8880,p8881);
FA fa2853(p8877,p8726,p8734,p8882,p8883);
HA ha1588(p8875,p8879,p8884,p8885);
FA fa2854(p8728,p8730,p8740,p8886,p8887);
FA fa2855(p8881,p8885,p8736,p8888,p8889);
HA ha1589(p8883,p8738,p8890,p8891);
FA fa2856(p8887,p8889,p8742,p8892,p8893);
FA fa2857(p8744,p8891,p8746,p8894,p8895);
HA ha1590(p8750,p8893,p8896,p8897);
FA fa2858(p8748,p8895,p8897,p8898,p8899);
HA ha1591(p8752,p8899,p8900,p8901);
FA fa2859(p8901,p8754,p8756,p8902,p8903);
FA fa2860(ip_19_63,ip_20_62,ip_21_61,p8904,p8905);
FA fa2861(ip_22_60,ip_23_59,ip_24_58,p8906,p8907);
FA fa2862(ip_25_57,ip_26_56,ip_27_55,p8908,p8909);
FA fa2863(ip_28_54,ip_29_53,ip_30_52,p8910,p8911);
FA fa2864(ip_31_51,ip_32_50,ip_33_49,p8912,p8913);
HA ha1592(ip_34_48,ip_35_47,p8914,p8915);
FA fa2865(ip_36_46,ip_37_45,ip_38_44,p8916,p8917);
FA fa2866(ip_39_43,ip_40_42,ip_41_41,p8918,p8919);
FA fa2867(ip_42_40,ip_43_39,ip_44_38,p8920,p8921);
FA fa2868(ip_45_37,ip_46_36,ip_47_35,p8922,p8923);
HA ha1593(ip_48_34,ip_49_33,p8924,p8925);
FA fa2869(ip_50_32,ip_51_31,ip_52_30,p8926,p8927);
FA fa2870(ip_53_29,ip_54_28,ip_55_27,p8928,p8929);
FA fa2871(ip_56_26,ip_57_25,ip_58_24,p8930,p8931);
HA ha1594(ip_59_23,ip_60_22,p8932,p8933);
FA fa2872(ip_61_21,ip_62_20,ip_63_19,p8934,p8935);
HA ha1595(p8766,p8772,p8936,p8937);
HA ha1596(p8774,p8776,p8938,p8939);
HA ha1597(p8778,p8780,p8940,p8941);
FA fa2873(p8788,p8790,p8794,p8942,p8943);
FA fa2874(p8915,p8925,p8933,p8944,p8945);
HA ha1598(p8802,p8804,p8946,p8947);
FA fa2875(p8905,p8907,p8909,p8948,p8949);
FA fa2876(p8911,p8913,p8917,p8950,p8951);
FA fa2877(p8919,p8921,p8923,p8952,p8953);
FA fa2878(p8927,p8929,p8931,p8954,p8955);
FA fa2879(p8935,p8937,p8939,p8956,p8957);
FA fa2880(p8941,p8760,p8762,p8958,p8959);
HA ha1599(p8764,p8768,p8960,p8961);
FA fa2881(p8770,p8782,p8784,p8962,p8963);
FA fa2882(p8786,p8792,p8814,p8964,p8965);
FA fa2883(p8943,p8945,p8947,p8966,p8967);
FA fa2884(p8796,p8798,p8800,p8968,p8969);
FA fa2885(p8806,p8949,p8951,p8970,p8971);
HA ha1600(p8953,p8955,p8972,p8973);
FA fa2886(p8957,p8961,p8808,p8974,p8975);
FA fa2887(p8810,p8812,p8816,p8976,p8977);
FA fa2888(p8834,p8836,p8959,p8978,p8979);
FA fa2889(p8963,p8965,p8967,p8980,p8981);
HA ha1601(p8973,p8818,p8982,p8983);
HA ha1602(p8820,p8822,p8984,p8985);
FA fa2890(p8824,p8826,p8828,p8986,p8987);
HA ha1603(p8830,p8844,p8988,p8989);
HA ha1604(p8846,p8969,p8990,p8991);
FA fa2891(p8971,p8975,p8832,p8992,p8993);
FA fa2892(p8838,p8850,p8977,p8994,p8995);
HA ha1605(p8979,p8981,p8996,p8997);
FA fa2893(p8983,p8985,p8989,p8998,p8999);
FA fa2894(p8991,p8840,p8842,p9000,p9001);
HA ha1606(p8848,p8862,p9002,p9003);
HA ha1607(p8987,p8993,p9004,p9005);
FA fa2895(p8997,p8852,p8854,p9006,p9007);
FA fa2896(p8856,p8858,p8995,p9008,p9009);
FA fa2897(p8999,p9003,p9005,p9010,p9011);
FA fa2898(p8860,p8872,p9001,p9012,p9013);
FA fa2899(p8864,p8866,p8868,p9014,p9015);
HA ha1608(p8876,p9007,p9016,p9017);
FA fa2900(p9009,p9011,p8870,p9018,p9019);
FA fa2901(p8878,p9013,p9017,p9020,p9021);
HA ha1609(p8874,p8884,p9022,p9023);
HA ha1610(p9015,p9019,p9024,p9025);
FA fa2902(p8880,p9021,p9023,p9026,p9027);
FA fa2903(p9025,p8882,p8886,p9028,p9029);
HA ha1611(p8888,p8890,p9030,p9031);
FA fa2904(p9027,p9029,p9031,p9032,p9033);
FA fa2905(p8892,p8896,p8894,p9034,p9035);
FA fa2906(p9033,p9035,p8898,p9036,p9037);
FA fa2907(p8900,p9037,p8902,p9038,p9039);
HA ha1612(ip_20_63,ip_21_62,p9040,p9041);
FA fa2908(ip_22_61,ip_23_60,ip_24_59,p9042,p9043);
FA fa2909(ip_25_58,ip_26_57,ip_27_56,p9044,p9045);
FA fa2910(ip_28_55,ip_29_54,ip_30_53,p9046,p9047);
FA fa2911(ip_31_52,ip_32_51,ip_33_50,p9048,p9049);
HA ha1613(ip_34_49,ip_35_48,p9050,p9051);
FA fa2912(ip_36_47,ip_37_46,ip_38_45,p9052,p9053);
FA fa2913(ip_39_44,ip_40_43,ip_41_42,p9054,p9055);
FA fa2914(ip_42_41,ip_43_40,ip_44_39,p9056,p9057);
FA fa2915(ip_45_38,ip_46_37,ip_47_36,p9058,p9059);
FA fa2916(ip_48_35,ip_49_34,ip_50_33,p9060,p9061);
FA fa2917(ip_51_32,ip_52_31,ip_53_30,p9062,p9063);
HA ha1614(ip_54_29,ip_55_28,p9064,p9065);
FA fa2918(ip_56_27,ip_57_26,ip_58_25,p9066,p9067);
HA ha1615(ip_59_24,ip_60_23,p9068,p9069);
FA fa2919(ip_61_22,ip_62_21,ip_63_20,p9070,p9071);
FA fa2920(p8914,p8924,p8932,p9072,p9073);
FA fa2921(p9041,p9051,p9065,p9074,p9075);
HA ha1616(p9069,p8936,p9076,p9077);
FA fa2922(p8938,p8940,p9043,p9078,p9079);
HA ha1617(p9045,p9047,p9080,p9081);
HA ha1618(p9049,p9053,p9082,p9083);
FA fa2923(p9055,p9057,p9059,p9084,p9085);
FA fa2924(p9061,p9063,p9067,p9086,p9087);
FA fa2925(p9071,p8904,p8906,p9088,p9089);
FA fa2926(p8908,p8910,p8912,p9090,p9091);
HA ha1619(p8916,p8918,p9092,p9093);
FA fa2927(p8920,p8922,p8926,p9094,p9095);
HA ha1620(p8928,p8930,p9096,p9097);
FA fa2928(p8934,p8946,p9073,p9098,p9099);
FA fa2929(p9075,p9077,p9081,p9100,p9101);
HA ha1621(p9083,p8942,p9102,p9103);
HA ha1622(p8944,p8960,p9104,p9105);
FA fa2930(p9079,p9085,p9087,p9106,p9107);
FA fa2931(p9093,p9097,p8948,p9108,p9109);
FA fa2932(p8950,p8952,p8954,p9110,p9111);
FA fa2933(p8956,p8972,p9089,p9112,p9113);
HA ha1623(p9091,p9095,p9114,p9115);
FA fa2934(p9099,p9101,p9103,p9116,p9117);
HA ha1624(p9105,p8958,p9118,p9119);
FA fa2935(p8962,p8964,p8966,p9120,p9121);
HA ha1625(p9107,p9109,p9122,p9123);
FA fa2936(p9115,p8968,p8970,p9124,p9125);
HA ha1626(p8974,p8982,p9126,p9127);
FA fa2937(p8984,p8988,p8990,p9128,p9129);
FA fa2938(p9111,p9113,p9117,p9130,p9131);
FA fa2939(p9119,p9123,p8976,p9132,p9133);
FA fa2940(p8978,p8980,p8996,p9134,p9135);
FA fa2941(p9121,p9127,p8986,p9136,p9137);
FA fa2942(p8992,p9002,p9004,p9138,p9139);
FA fa2943(p9125,p9129,p9131,p9140,p9141);
HA ha1627(p9133,p8994,p9142,p9143);
FA fa2944(p8998,p9135,p9137,p9144,p9145);
FA fa2945(p9000,p9139,p9141,p9146,p9147);
FA fa2946(p9143,p9006,p9008,p9148,p9149);
FA fa2947(p9010,p9016,p9145,p9150,p9151);
FA fa2948(p9012,p9147,p9014,p9152,p9153);
HA ha1628(p9018,p9022,p9154,p9155);
FA fa2949(p9024,p9149,p9151,p9156,p9157);
HA ha1629(p9020,p9153,p9158,p9159);
HA ha1630(p9155,p9157,p9160,p9161);
FA fa2950(p9159,p9026,p9030,p9162,p9163);
FA fa2951(p9161,p9028,p9163,p9164,p9165);
FA fa2952(p9032,p9165,p9034,p9166,p9167);
FA fa2953(p9167,p9036,p9038,p9168,p9169);
HA ha1631(ip_21_63,ip_22_62,p9170,p9171);
FA fa2954(ip_23_61,ip_24_60,ip_25_59,p9172,p9173);
FA fa2955(ip_26_58,ip_27_57,ip_28_56,p9174,p9175);
FA fa2956(ip_29_55,ip_30_54,ip_31_53,p9176,p9177);
HA ha1632(ip_32_52,ip_33_51,p9178,p9179);
HA ha1633(ip_34_50,ip_35_49,p9180,p9181);
HA ha1634(ip_36_48,ip_37_47,p9182,p9183);
HA ha1635(ip_38_46,ip_39_45,p9184,p9185);
HA ha1636(ip_40_44,ip_41_43,p9186,p9187);
FA fa2957(ip_42_42,ip_43_41,ip_44_40,p9188,p9189);
HA ha1637(ip_45_39,ip_46_38,p9190,p9191);
HA ha1638(ip_47_37,ip_48_36,p9192,p9193);
FA fa2958(ip_49_35,ip_50_34,ip_51_33,p9194,p9195);
FA fa2959(ip_52_32,ip_53_31,ip_54_30,p9196,p9197);
HA ha1639(ip_55_29,ip_56_28,p9198,p9199);
FA fa2960(ip_57_27,ip_58_26,ip_59_25,p9200,p9201);
FA fa2961(ip_60_24,ip_61_23,ip_62_22,p9202,p9203);
HA ha1640(ip_63_21,p9040,p9204,p9205);
HA ha1641(p9050,p9064,p9206,p9207);
HA ha1642(p9068,p9171,p9208,p9209);
HA ha1643(p9179,p9181,p9210,p9211);
FA fa2962(p9183,p9185,p9187,p9212,p9213);
FA fa2963(p9191,p9193,p9199,p9214,p9215);
FA fa2964(p9173,p9175,p9177,p9216,p9217);
FA fa2965(p9189,p9195,p9197,p9218,p9219);
HA ha1644(p9201,p9203,p9220,p9221);
FA fa2966(p9205,p9207,p9209,p9222,p9223);
FA fa2967(p9211,p9042,p9044,p9224,p9225);
FA fa2968(p9046,p9048,p9052,p9226,p9227);
FA fa2969(p9054,p9056,p9058,p9228,p9229);
FA fa2970(p9060,p9062,p9066,p9230,p9231);
FA fa2971(p9070,p9076,p9080,p9232,p9233);
FA fa2972(p9082,p9213,p9215,p9234,p9235);
FA fa2973(p9221,p9072,p9074,p9236,p9237);
FA fa2974(p9092,p9096,p9217,p9238,p9239);
FA fa2975(p9219,p9223,p9078,p9240,p9241);
HA ha1645(p9084,p9086,p9242,p9243);
FA fa2976(p9102,p9104,p9225,p9244,p9245);
FA fa2977(p9227,p9229,p9231,p9246,p9247);
HA ha1646(p9233,p9235,p9248,p9249);
FA fa2978(p9088,p9090,p9094,p9250,p9251);
HA ha1647(p9098,p9100,p9252,p9253);
FA fa2979(p9114,p9237,p9239,p9254,p9255);
FA fa2980(p9241,p9243,p9249,p9256,p9257);
FA fa2981(p9106,p9108,p9118,p9258,p9259);
HA ha1648(p9122,p9245,p9260,p9261);
FA fa2982(p9247,p9253,p9110,p9262,p9263);
HA ha1649(p9112,p9116,p9264,p9265);
FA fa2983(p9126,p9251,p9255,p9266,p9267);
FA fa2984(p9257,p9261,p9120,p9268,p9269);
HA ha1650(p9259,p9263,p9270,p9271);
HA ha1651(p9265,p9124,p9272,p9273);
FA fa2985(p9128,p9130,p9132,p9274,p9275);
HA ha1652(p9267,p9269,p9276,p9277);
HA ha1653(p9271,p9134,p9278,p9279);
FA fa2986(p9136,p9142,p9273,p9280,p9281);
FA fa2987(p9277,p9138,p9140,p9282,p9283);
FA fa2988(p9275,p9279,p9144,p9284,p9285);
HA ha1654(p9281,p9146,p9286,p9287);
FA fa2989(p9283,p9285,p9148,p9288,p9289);
FA fa2990(p9150,p9154,p9287,p9290,p9291);
FA fa2991(p9152,p9158,p9289,p9292,p9293);
HA ha1655(p9156,p9160,p9294,p9295);
FA fa2992(p9291,p9293,p9295,p9296,p9297);
HA ha1656(p9162,p9297,p9298,p9299);
HA ha1657(p9164,p9299,p9300,p9301);
FA fa2993(p9301,p9166,p9168,p9302,p9303);
HA ha1658(ip_22_63,ip_23_62,p9304,p9305);
FA fa2994(ip_24_61,ip_25_60,ip_26_59,p9306,p9307);
HA ha1659(ip_27_58,ip_28_57,p9308,p9309);
HA ha1660(ip_29_56,ip_30_55,p9310,p9311);
FA fa2995(ip_31_54,ip_32_53,ip_33_52,p9312,p9313);
FA fa2996(ip_34_51,ip_35_50,ip_36_49,p9314,p9315);
FA fa2997(ip_37_48,ip_38_47,ip_39_46,p9316,p9317);
FA fa2998(ip_40_45,ip_41_44,ip_42_43,p9318,p9319);
FA fa2999(ip_43_42,ip_44_41,ip_45_40,p9320,p9321);
FA fa3000(ip_46_39,ip_47_38,ip_48_37,p9322,p9323);
FA fa3001(ip_49_36,ip_50_35,ip_51_34,p9324,p9325);
FA fa3002(ip_52_33,ip_53_32,ip_54_31,p9326,p9327);
HA ha1661(ip_55_30,ip_56_29,p9328,p9329);
HA ha1662(ip_57_28,ip_58_27,p9330,p9331);
FA fa3003(ip_59_26,ip_60_25,ip_61_24,p9332,p9333);
FA fa3004(ip_62_23,ip_63_22,p9170,p9334,p9335);
FA fa3005(p9178,p9180,p9182,p9336,p9337);
FA fa3006(p9184,p9186,p9190,p9338,p9339);
FA fa3007(p9192,p9198,p9305,p9340,p9341);
HA ha1663(p9309,p9311,p9342,p9343);
FA fa3008(p9329,p9331,p9204,p9344,p9345);
FA fa3009(p9206,p9208,p9210,p9346,p9347);
FA fa3010(p9307,p9313,p9315,p9348,p9349);
FA fa3011(p9317,p9319,p9321,p9350,p9351);
HA ha1664(p9323,p9325,p9352,p9353);
FA fa3012(p9327,p9333,p9335,p9354,p9355);
HA ha1665(p9343,p9172,p9356,p9357);
FA fa3013(p9174,p9176,p9188,p9358,p9359);
FA fa3014(p9194,p9196,p9200,p9360,p9361);
HA ha1666(p9202,p9220,p9362,p9363);
HA ha1667(p9337,p9339,p9364,p9365);
FA fa3015(p9341,p9345,p9353,p9366,p9367);
HA ha1668(p9212,p9214,p9368,p9369);
HA ha1669(p9347,p9349,p9370,p9371);
FA fa3016(p9351,p9355,p9357,p9372,p9373);
FA fa3017(p9363,p9365,p9216,p9374,p9375);
HA ha1670(p9218,p9222,p9376,p9377);
FA fa3018(p9359,p9361,p9367,p9378,p9379);
FA fa3019(p9369,p9371,p9224,p9380,p9381);
FA fa3020(p9226,p9228,p9230,p9382,p9383);
FA fa3021(p9232,p9234,p9242,p9384,p9385);
HA ha1671(p9248,p9373,p9386,p9387);
FA fa3022(p9375,p9377,p9236,p9388,p9389);
FA fa3023(p9238,p9240,p9252,p9390,p9391);
FA fa3024(p9379,p9381,p9387,p9392,p9393);
FA fa3025(p9244,p9246,p9260,p9394,p9395);
FA fa3026(p9383,p9385,p9389,p9396,p9397);
FA fa3027(p9250,p9254,p9256,p9398,p9399);
HA ha1672(p9264,p9391,p9400,p9401);
FA fa3028(p9393,p9258,p9262,p9402,p9403);
FA fa3029(p9270,p9395,p9397,p9404,p9405);
FA fa3030(p9401,p9266,p9268,p9406,p9407);
HA ha1673(p9272,p9276,p9408,p9409);
HA ha1674(p9399,p9278,p9410,p9411);
FA fa3031(p9403,p9405,p9409,p9412,p9413);
FA fa3032(p9274,p9407,p9411,p9414,p9415);
FA fa3033(p9280,p9413,p9282,p9416,p9417);
FA fa3034(p9284,p9286,p9415,p9418,p9419);
HA ha1675(p9417,p9288,p9420,p9421);
FA fa3035(p9419,p9290,p9294,p9422,p9423);
HA ha1676(p9421,p9292,p9424,p9425);
HA ha1677(p9423,p9425,p9426,p9427);
FA fa3036(p9296,p9298,p9427,p9428,p9429);
FA fa3037(p9300,p9429,p9302,p9430,p9431);
HA ha1678(ip_23_63,ip_24_62,p9432,p9433);
FA fa3038(ip_25_61,ip_26_60,ip_27_59,p9434,p9435);
HA ha1679(ip_28_58,ip_29_57,p9436,p9437);
FA fa3039(ip_30_56,ip_31_55,ip_32_54,p9438,p9439);
HA ha1680(ip_33_53,ip_34_52,p9440,p9441);
FA fa3040(ip_35_51,ip_36_50,ip_37_49,p9442,p9443);
FA fa3041(ip_38_48,ip_39_47,ip_40_46,p9444,p9445);
HA ha1681(ip_41_45,ip_42_44,p9446,p9447);
FA fa3042(ip_43_43,ip_44_42,ip_45_41,p9448,p9449);
FA fa3043(ip_46_40,ip_47_39,ip_48_38,p9450,p9451);
HA ha1682(ip_49_37,ip_50_36,p9452,p9453);
HA ha1683(ip_51_35,ip_52_34,p9454,p9455);
FA fa3044(ip_53_33,ip_54_32,ip_55_31,p9456,p9457);
FA fa3045(ip_56_30,ip_57_29,ip_58_28,p9458,p9459);
FA fa3046(ip_59_27,ip_60_26,ip_61_25,p9460,p9461);
FA fa3047(ip_62_24,ip_63_23,p9304,p9462,p9463);
FA fa3048(p9308,p9310,p9328,p9464,p9465);
HA ha1684(p9330,p9433,p9466,p9467);
HA ha1685(p9437,p9441,p9468,p9469);
HA ha1686(p9447,p9453,p9470,p9471);
HA ha1687(p9455,p9342,p9472,p9473);
FA fa3049(p9435,p9439,p9443,p9474,p9475);
FA fa3050(p9445,p9449,p9451,p9476,p9477);
FA fa3051(p9457,p9459,p9461,p9478,p9479);
FA fa3052(p9463,p9467,p9469,p9480,p9481);
HA ha1688(p9471,p9306,p9482,p9483);
FA fa3053(p9312,p9314,p9316,p9484,p9485);
FA fa3054(p9318,p9320,p9322,p9486,p9487);
FA fa3055(p9324,p9326,p9332,p9488,p9489);
FA fa3056(p9334,p9352,p9465,p9490,p9491);
FA fa3057(p9473,p9336,p9338,p9492,p9493);
FA fa3058(p9340,p9344,p9356,p9494,p9495);
FA fa3059(p9362,p9364,p9475,p9496,p9497);
HA ha1689(p9477,p9479,p9498,p9499);
FA fa3060(p9481,p9483,p9346,p9500,p9501);
FA fa3061(p9348,p9350,p9354,p9502,p9503);
FA fa3062(p9368,p9370,p9485,p9504,p9505);
FA fa3063(p9487,p9489,p9491,p9506,p9507);
HA ha1690(p9499,p9358,p9508,p9509);
FA fa3064(p9360,p9366,p9376,p9510,p9511);
FA fa3065(p9493,p9495,p9497,p9512,p9513);
FA fa3066(p9501,p9372,p9374,p9514,p9515);
HA ha1691(p9386,p9503,p9516,p9517);
HA ha1692(p9505,p9507,p9518,p9519);
FA fa3067(p9509,p9378,p9380,p9520,p9521);
FA fa3068(p9511,p9513,p9517,p9522,p9523);
HA ha1693(p9519,p9382,p9524,p9525);
FA fa3069(p9384,p9388,p9515,p9526,p9527);
FA fa3070(p9390,p9392,p9400,p9528,p9529);
HA ha1694(p9521,p9523,p9530,p9531);
FA fa3071(p9525,p9394,p9396,p9532,p9533);
FA fa3072(p9527,p9531,p9398,p9534,p9535);
HA ha1695(p9408,p9529,p9536,p9537);
HA ha1696(p9402,p9404,p9538,p9539);
HA ha1697(p9410,p9533,p9540,p9541);
FA fa3073(p9535,p9537,p9406,p9542,p9543);
FA fa3074(p9539,p9541,p9412,p9544,p9545);
HA ha1698(p9543,p9414,p9546,p9547);
FA fa3075(p9545,p9416,p9547,p9548,p9549);
HA ha1699(p9418,p9420,p9550,p9551);
FA fa3076(p9549,p9551,p9424,p9552,p9553);
FA fa3077(p9422,p9426,p9553,p9554,p9555);
FA fa3078(p9555,p9428,p9430,p9556,p9557);
FA fa3079(ip_24_63,ip_25_62,ip_26_61,p9558,p9559);
HA ha1700(ip_27_60,ip_28_59,p9560,p9561);
HA ha1701(ip_29_58,ip_30_57,p9562,p9563);
FA fa3080(ip_31_56,ip_32_55,ip_33_54,p9564,p9565);
HA ha1702(ip_34_53,ip_35_52,p9566,p9567);
HA ha1703(ip_36_51,ip_37_50,p9568,p9569);
FA fa3081(ip_38_49,ip_39_48,ip_40_47,p9570,p9571);
HA ha1704(ip_41_46,ip_42_45,p9572,p9573);
FA fa3082(ip_43_44,ip_44_43,ip_45_42,p9574,p9575);
HA ha1705(ip_46_41,ip_47_40,p9576,p9577);
FA fa3083(ip_48_39,ip_49_38,ip_50_37,p9578,p9579);
HA ha1706(ip_51_36,ip_52_35,p9580,p9581);
FA fa3084(ip_53_34,ip_54_33,ip_55_32,p9582,p9583);
FA fa3085(ip_56_31,ip_57_30,ip_58_29,p9584,p9585);
FA fa3086(ip_59_28,ip_60_27,ip_61_26,p9586,p9587);
FA fa3087(ip_62_25,ip_63_24,p9432,p9588,p9589);
FA fa3088(p9436,p9440,p9446,p9590,p9591);
HA ha1707(p9452,p9454,p9592,p9593);
HA ha1708(p9561,p9563,p9594,p9595);
FA fa3089(p9567,p9569,p9573,p9596,p9597);
HA ha1709(p9577,p9581,p9598,p9599);
HA ha1710(p9466,p9468,p9600,p9601);
HA ha1711(p9470,p9559,p9602,p9603);
FA fa3090(p9565,p9571,p9575,p9604,p9605);
HA ha1712(p9579,p9583,p9606,p9607);
FA fa3091(p9585,p9587,p9589,p9608,p9609);
HA ha1713(p9593,p9595,p9610,p9611);
HA ha1714(p9599,p9434,p9612,p9613);
HA ha1715(p9438,p9442,p9614,p9615);
FA fa3092(p9444,p9448,p9450,p9616,p9617);
HA ha1716(p9456,p9458,p9618,p9619);
FA fa3093(p9460,p9462,p9472,p9620,p9621);
FA fa3094(p9591,p9597,p9601,p9622,p9623);
HA ha1717(p9603,p9607,p9624,p9625);
FA fa3095(p9611,p9464,p9482,p9626,p9627);
FA fa3096(p9605,p9609,p9613,p9628,p9629);
FA fa3097(p9615,p9619,p9625,p9630,p9631);
FA fa3098(p9474,p9476,p9478,p9632,p9633);
HA ha1718(p9480,p9498,p9634,p9635);
FA fa3099(p9617,p9621,p9623,p9636,p9637);
FA fa3100(p9484,p9486,p9488,p9638,p9639);
HA ha1719(p9490,p9627,p9640,p9641);
HA ha1720(p9629,p9631,p9642,p9643);
HA ha1721(p9635,p9492,p9644,p9645);
FA fa3101(p9494,p9496,p9500,p9646,p9647);
HA ha1722(p9508,p9633,p9648,p9649);
FA fa3102(p9637,p9641,p9643,p9650,p9651);
FA fa3103(p9502,p9504,p9506,p9652,p9653);
FA fa3104(p9516,p9518,p9639,p9654,p9655);
HA ha1723(p9645,p9649,p9656,p9657);
HA ha1724(p9510,p9512,p9658,p9659);
HA ha1725(p9647,p9651,p9660,p9661);
FA fa3105(p9657,p9514,p9524,p9662,p9663);
FA fa3106(p9653,p9655,p9659,p9664,p9665);
FA fa3107(p9661,p9520,p9522,p9666,p9667);
FA fa3108(p9530,p9526,p9663,p9668,p9669);
FA fa3109(p9665,p9528,p9536,p9670,p9671);
HA ha1726(p9667,p9532,p9672,p9673);
HA ha1727(p9534,p9538,p9674,p9675);
FA fa3110(p9540,p9669,p9671,p9676,p9677);
HA ha1728(p9673,p9675,p9678,p9679);
HA ha1729(p9542,p9677,p9680,p9681);
HA ha1730(p9679,p9544,p9682,p9683);
HA ha1731(p9546,p9681,p9684,p9685);
HA ha1732(p9683,p9685,p9686,p9687);
FA fa3111(p9550,p9687,p9548,p9688,p9689);
FA fa3112(p9689,p9552,p9554,p9690,p9691);
FA fa3113(ip_25_63,ip_26_62,ip_27_61,p9692,p9693);
HA ha1733(ip_28_60,ip_29_59,p9694,p9695);
HA ha1734(ip_30_58,ip_31_57,p9696,p9697);
HA ha1735(ip_32_56,ip_33_55,p9698,p9699);
HA ha1736(ip_34_54,ip_35_53,p9700,p9701);
FA fa3114(ip_36_52,ip_37_51,ip_38_50,p9702,p9703);
FA fa3115(ip_39_49,ip_40_48,ip_41_47,p9704,p9705);
FA fa3116(ip_42_46,ip_43_45,ip_44_44,p9706,p9707);
HA ha1737(ip_45_43,ip_46_42,p9708,p9709);
HA ha1738(ip_47_41,ip_48_40,p9710,p9711);
FA fa3117(ip_49_39,ip_50_38,ip_51_37,p9712,p9713);
HA ha1739(ip_52_36,ip_53_35,p9714,p9715);
HA ha1740(ip_54_34,ip_55_33,p9716,p9717);
HA ha1741(ip_56_32,ip_57_31,p9718,p9719);
HA ha1742(ip_58_30,ip_59_29,p9720,p9721);
HA ha1743(ip_60_28,ip_61_27,p9722,p9723);
HA ha1744(ip_62_26,ip_63_25,p9724,p9725);
FA fa3118(p9560,p9562,p9566,p9726,p9727);
FA fa3119(p9568,p9572,p9576,p9728,p9729);
FA fa3120(p9580,p9695,p9697,p9730,p9731);
HA ha1745(p9699,p9701,p9732,p9733);
HA ha1746(p9709,p9711,p9734,p9735);
FA fa3121(p9715,p9717,p9719,p9736,p9737);
FA fa3122(p9721,p9723,p9725,p9738,p9739);
FA fa3123(p9592,p9594,p9598,p9740,p9741);
FA fa3124(p9693,p9703,p9705,p9742,p9743);
HA ha1747(p9707,p9713,p9744,p9745);
FA fa3125(p9733,p9735,p9558,p9746,p9747);
HA ha1748(p9564,p9570,p9748,p9749);
FA fa3126(p9574,p9578,p9582,p9750,p9751);
FA fa3127(p9584,p9586,p9588,p9752,p9753);
FA fa3128(p9600,p9602,p9606,p9754,p9755);
FA fa3129(p9610,p9727,p9729,p9756,p9757);
FA fa3130(p9731,p9737,p9739,p9758,p9759);
FA fa3131(p9745,p9590,p9596,p9760,p9761);
FA fa3132(p9612,p9614,p9618,p9762,p9763);
FA fa3133(p9624,p9741,p9743,p9764,p9765);
HA ha1749(p9747,p9749,p9766,p9767);
FA fa3134(p9604,p9608,p9751,p9768,p9769);
FA fa3135(p9753,p9755,p9757,p9770,p9771);
FA fa3136(p9759,p9767,p9616,p9772,p9773);
HA ha1750(p9620,p9622,p9774,p9775);
HA ha1751(p9634,p9761,p9776,p9777);
HA ha1752(p9763,p9765,p9778,p9779);
HA ha1753(p9626,p9628,p9780,p9781);
FA fa3137(p9630,p9640,p9642,p9782,p9783);
FA fa3138(p9769,p9771,p9773,p9784,p9785);
FA fa3139(p9775,p9777,p9779,p9786,p9787);
FA fa3140(p9632,p9636,p9644,p9788,p9789);
FA fa3141(p9648,p9781,p9638,p9790,p9791);
FA fa3142(p9656,p9783,p9785,p9792,p9793);
FA fa3143(p9787,p9646,p9650,p9794,p9795);
FA fa3144(p9658,p9660,p9789,p9796,p9797);
FA fa3145(p9791,p9652,p9654,p9798,p9799);
FA fa3146(p9793,p9795,p9797,p9800,p9801);
FA fa3147(p9662,p9664,p9799,p9802,p9803);
FA fa3148(p9666,p9801,p9668,p9804,p9805);
FA fa3149(p9672,p9674,p9803,p9806,p9807);
HA ha1754(p9670,p9678,p9808,p9809);
HA ha1755(p9805,p9676,p9810,p9811);
HA ha1756(p9680,p9807,p9812,p9813);
FA fa3150(p9809,p9682,p9684,p9814,p9815);
FA fa3151(p9811,p9813,p9686,p9816,p9817);
FA fa3152(p9815,p9817,p9688,p9818,p9819);
HA ha1757(ip_26_63,ip_27_62,p9820,p9821);
FA fa3153(ip_28_61,ip_29_60,ip_30_59,p9822,p9823);
HA ha1758(ip_31_58,ip_32_57,p9824,p9825);
FA fa3154(ip_33_56,ip_34_55,ip_35_54,p9826,p9827);
FA fa3155(ip_36_53,ip_37_52,ip_38_51,p9828,p9829);
FA fa3156(ip_39_50,ip_40_49,ip_41_48,p9830,p9831);
FA fa3157(ip_42_47,ip_43_46,ip_44_45,p9832,p9833);
FA fa3158(ip_45_44,ip_46_43,ip_47_42,p9834,p9835);
FA fa3159(ip_48_41,ip_49_40,ip_50_39,p9836,p9837);
FA fa3160(ip_51_38,ip_52_37,ip_53_36,p9838,p9839);
FA fa3161(ip_54_35,ip_55_34,ip_56_33,p9840,p9841);
FA fa3162(ip_57_32,ip_58_31,ip_59_30,p9842,p9843);
FA fa3163(ip_60_29,ip_61_28,ip_62_27,p9844,p9845);
HA ha1759(ip_63_26,p9694,p9846,p9847);
HA ha1760(p9696,p9698,p9848,p9849);
HA ha1761(p9700,p9708,p9850,p9851);
FA fa3164(p9710,p9714,p9716,p9852,p9853);
FA fa3165(p9718,p9720,p9722,p9854,p9855);
FA fa3166(p9724,p9821,p9825,p9856,p9857);
FA fa3167(p9732,p9734,p9823,p9858,p9859);
FA fa3168(p9827,p9829,p9831,p9860,p9861);
FA fa3169(p9833,p9835,p9837,p9862,p9863);
FA fa3170(p9839,p9841,p9843,p9864,p9865);
FA fa3171(p9845,p9847,p9849,p9866,p9867);
FA fa3172(p9851,p9692,p9702,p9868,p9869);
FA fa3173(p9704,p9706,p9712,p9870,p9871);
FA fa3174(p9744,p9853,p9855,p9872,p9873);
HA ha1762(p9857,p9726,p9874,p9875);
HA ha1763(p9728,p9730,p9876,p9877);
FA fa3175(p9736,p9738,p9748,p9878,p9879);
FA fa3176(p9859,p9861,p9863,p9880,p9881);
HA ha1764(p9865,p9867,p9882,p9883);
FA fa3177(p9740,p9742,p9746,p9884,p9885);
FA fa3178(p9766,p9869,p9871,p9886,p9887);
FA fa3179(p9873,p9875,p9877,p9888,p9889);
FA fa3180(p9883,p9750,p9752,p9890,p9891);
FA fa3181(p9754,p9756,p9758,p9892,p9893);
FA fa3182(p9879,p9881,p9760,p9894,p9895);
HA ha1765(p9762,p9764,p9896,p9897);
FA fa3183(p9774,p9776,p9778,p9898,p9899);
FA fa3184(p9885,p9887,p9889,p9900,p9901);
HA ha1766(p9768,p9770,p9902,p9903);
FA fa3185(p9772,p9780,p9891,p9904,p9905);
HA ha1767(p9893,p9895,p9906,p9907);
HA ha1768(p9897,p9899,p9908,p9909);
FA fa3186(p9901,p9903,p9907,p9910,p9911);
FA fa3187(p9782,p9784,p9786,p9912,p9913);
FA fa3188(p9905,p9909,p9788,p9914,p9915);
HA ha1769(p9790,p9911,p9916,p9917);
HA ha1770(p9792,p9913,p9918,p9919);
HA ha1771(p9915,p9917,p9920,p9921);
FA fa3189(p9794,p9796,p9919,p9922,p9923);
FA fa3190(p9921,p9798,p9800,p9924,p9925);
HA ha1772(p9923,p9802,p9926,p9927);
FA fa3191(p9925,p9804,p9808,p9928,p9929);
FA fa3192(p9927,p9806,p9810,p9930,p9931);
FA fa3193(p9812,p9929,p9931,p9932,p9933);
HA ha1773(p9814,p9816,p9934,p9935);
FA fa3194(p9933,p9935,p9818,p9936,p9937);
FA fa3195(ip_27_63,ip_28_62,ip_29_61,p9938,p9939);
FA fa3196(ip_30_60,ip_31_59,ip_32_58,p9940,p9941);
FA fa3197(ip_33_57,ip_34_56,ip_35_55,p9942,p9943);
FA fa3198(ip_36_54,ip_37_53,ip_38_52,p9944,p9945);
FA fa3199(ip_39_51,ip_40_50,ip_41_49,p9946,p9947);
FA fa3200(ip_42_48,ip_43_47,ip_44_46,p9948,p9949);
FA fa3201(ip_45_45,ip_46_44,ip_47_43,p9950,p9951);
HA ha1774(ip_48_42,ip_49_41,p9952,p9953);
HA ha1775(ip_50_40,ip_51_39,p9954,p9955);
FA fa3202(ip_52_38,ip_53_37,ip_54_36,p9956,p9957);
FA fa3203(ip_55_35,ip_56_34,ip_57_33,p9958,p9959);
HA ha1776(ip_58_32,ip_59_31,p9960,p9961);
FA fa3204(ip_60_30,ip_61_29,ip_62_28,p9962,p9963);
FA fa3205(ip_63_27,p9820,p9824,p9964,p9965);
HA ha1777(p9953,p9955,p9966,p9967);
HA ha1778(p9961,p9846,p9968,p9969);
FA fa3206(p9848,p9850,p9939,p9970,p9971);
FA fa3207(p9941,p9943,p9945,p9972,p9973);
FA fa3208(p9947,p9949,p9951,p9974,p9975);
FA fa3209(p9957,p9959,p9963,p9976,p9977);
FA fa3210(p9967,p9822,p9826,p9978,p9979);
HA ha1779(p9828,p9830,p9980,p9981);
FA fa3211(p9832,p9834,p9836,p9982,p9983);
FA fa3212(p9838,p9840,p9842,p9984,p9985);
HA ha1780(p9844,p9965,p9986,p9987);
HA ha1781(p9969,p9852,p9988,p9989);
HA ha1782(p9854,p9856,p9990,p9991);
FA fa3213(p9971,p9973,p9975,p9992,p9993);
HA ha1783(p9977,p9981,p9994,p9995);
FA fa3214(p9987,p9858,p9860,p9996,p9997);
FA fa3215(p9862,p9864,p9866,p9998,p9999);
FA fa3216(p9874,p9876,p9882,p10000,p10001);
HA ha1784(p9979,p9983,p10002,p10003);
HA ha1785(p9985,p9989,p10004,p10005);
HA ha1786(p9991,p9995,p10006,p10007);
HA ha1787(p10003,p10005,p10008,p10009);
HA ha1788(p10007,p9868,p10010,p10011);
HA ha1789(p9870,p9872,p10012,p10013);
FA fa3217(p9993,p10001,p10009,p10014,p10015);
FA fa3218(p10011,p10013,p9878,p10016,p10017);
FA fa3219(p9880,p9997,p9999,p10018,p10019);
HA ha1790(p9884,p9886,p10020,p10021);
FA fa3220(p9888,p9896,p10015,p10022,p10023);
FA fa3221(p10017,p10019,p10021,p10024,p10025);
HA ha1791(p9890,p9892,p10026,p10027);
HA ha1792(p9894,p9902,p10028,p10029);
FA fa3222(p9906,p10023,p10027,p10030,p10031);
HA ha1793(p10029,p9898,p10032,p10033);
HA ha1794(p9900,p9908,p10034,p10035);
FA fa3223(p10025,p10033,p10035,p10036,p10037);
FA fa3224(p9904,p10031,p9910,p10038,p10039);
HA ha1795(p9916,p10037,p10040,p10041);
FA fa3225(p9912,p9914,p9918,p10042,p10043);
FA fa3226(p9920,p10039,p10041,p10044,p10045);
HA ha1796(p10043,p10045,p10046,p10047);
FA fa3227(p9922,p10047,p9924,p10048,p10049);
FA fa3228(p9926,p10049,p9928,p10050,p10051);
HA ha1797(p10051,p9930,p10052,p10053);
HA ha1798(p10053,p9932,p10054,p10055);
FA fa3229(p9934,p10055,p9936,p10056,p10057);
HA ha1799(ip_28_63,ip_29_62,p10058,p10059);
FA fa3230(ip_30_61,ip_31_60,ip_32_59,p10060,p10061);
FA fa3231(ip_33_58,ip_34_57,ip_35_56,p10062,p10063);
FA fa3232(ip_36_55,ip_37_54,ip_38_53,p10064,p10065);
FA fa3233(ip_39_52,ip_40_51,ip_41_50,p10066,p10067);
HA ha1800(ip_42_49,ip_43_48,p10068,p10069);
HA ha1801(ip_44_47,ip_45_46,p10070,p10071);
FA fa3234(ip_46_45,ip_47_44,ip_48_43,p10072,p10073);
FA fa3235(ip_49_42,ip_50_41,ip_51_40,p10074,p10075);
FA fa3236(ip_52_39,ip_53_38,ip_54_37,p10076,p10077);
HA ha1802(ip_55_36,ip_56_35,p10078,p10079);
HA ha1803(ip_57_34,ip_58_33,p10080,p10081);
FA fa3237(ip_59_32,ip_60_31,ip_61_30,p10082,p10083);
HA ha1804(ip_62_29,ip_63_28,p10084,p10085);
FA fa3238(p10059,p10069,p10071,p10086,p10087);
FA fa3239(p10079,p10081,p10085,p10088,p10089);
FA fa3240(p9952,p9954,p9960,p10090,p10091);
FA fa3241(p10061,p10063,p10065,p10092,p10093);
FA fa3242(p10067,p10073,p10075,p10094,p10095);
FA fa3243(p10077,p10083,p9966,p10096,p10097);
HA ha1805(p10087,p10089,p10098,p10099);
FA fa3244(p10091,p9938,p9940,p10100,p10101);
HA ha1806(p9942,p9944,p10102,p10103);
FA fa3245(p9946,p9948,p9950,p10104,p10105);
HA ha1807(p9956,p9958,p10106,p10107);
FA fa3246(p9962,p9968,p10093,p10108,p10109);
FA fa3247(p10095,p10097,p10099,p10110,p10111);
FA fa3248(p10103,p10107,p9964,p10112,p10113);
FA fa3249(p9980,p9986,p10101,p10114,p10115);
HA ha1808(p10105,p10109,p10116,p10117);
FA fa3250(p9970,p9972,p9974,p10118,p10119);
FA fa3251(p9976,p9988,p9990,p10120,p10121);
FA fa3252(p9994,p10002,p10004,p10122,p10123);
FA fa3253(p10006,p10111,p10113,p10124,p10125);
FA fa3254(p10115,p10117,p9978,p10126,p10127);
FA fa3255(p9982,p9984,p10008,p10128,p10129);
HA ha1809(p10010,p10012,p10130,p10131);
FA fa3256(p10119,p10121,p9992,p10132,p10133);
FA fa3257(p10000,p10123,p10125,p10134,p10135);
FA fa3258(p10127,p10129,p10131,p10136,p10137);
FA fa3259(p9996,p9998,p10020,p10138,p10139);
FA fa3260(p10133,p10014,p10016,p10140,p10141);
HA ha1810(p10018,p10026,p10142,p10143);
FA fa3261(p10028,p10135,p10137,p10144,p10145);
HA ha1811(p10139,p10022,p10146,p10147);
FA fa3262(p10032,p10034,p10143,p10148,p10149);
FA fa3263(p10024,p10141,p10145,p10150,p10151);
FA fa3264(p10147,p10030,p10149,p10152,p10153);
FA fa3265(p10036,p10040,p10151,p10154,p10155);
HA ha1812(p10038,p10153,p10156,p10157);
FA fa3266(p10042,p10155,p10157,p10158,p10159);
FA fa3267(p10044,p10046,p10159,p10160,p10161);
FA fa3268(p10161,p10048,p10050,p10162,p10163);
FA fa3269(p10052,p10054,p10163,p10164,p10165);
FA fa3270(ip_29_63,ip_30_62,ip_31_61,p10166,p10167);
FA fa3271(ip_32_60,ip_33_59,ip_34_58,p10168,p10169);
HA ha1813(ip_35_57,ip_36_56,p10170,p10171);
HA ha1814(ip_37_55,ip_38_54,p10172,p10173);
FA fa3272(ip_39_53,ip_40_52,ip_41_51,p10174,p10175);
FA fa3273(ip_42_50,ip_43_49,ip_44_48,p10176,p10177);
HA ha1815(ip_45_47,ip_46_46,p10178,p10179);
FA fa3274(ip_47_45,ip_48_44,ip_49_43,p10180,p10181);
HA ha1816(ip_50_42,ip_51_41,p10182,p10183);
HA ha1817(ip_52_40,ip_53_39,p10184,p10185);
FA fa3275(ip_54_38,ip_55_37,ip_56_36,p10186,p10187);
FA fa3276(ip_57_35,ip_58_34,ip_59_33,p10188,p10189);
FA fa3277(ip_60_32,ip_61_31,ip_62_30,p10190,p10191);
FA fa3278(ip_63_29,p10058,p10068,p10192,p10193);
FA fa3279(p10070,p10078,p10080,p10194,p10195);
HA ha1818(p10084,p10171,p10196,p10197);
HA ha1819(p10173,p10179,p10198,p10199);
FA fa3280(p10183,p10185,p10167,p10200,p10201);
HA ha1820(p10169,p10175,p10202,p10203);
HA ha1821(p10177,p10181,p10204,p10205);
HA ha1822(p10187,p10189,p10206,p10207);
HA ha1823(p10191,p10197,p10208,p10209);
FA fa3281(p10199,p10060,p10062,p10210,p10211);
HA ha1824(p10064,p10066,p10212,p10213);
FA fa3282(p10072,p10074,p10076,p10214,p10215);
FA fa3283(p10082,p10193,p10195,p10216,p10217);
FA fa3284(p10201,p10203,p10205,p10218,p10219);
FA fa3285(p10207,p10209,p10086,p10220,p10221);
HA ha1825(p10088,p10090,p10222,p10223);
HA ha1826(p10098,p10102,p10224,p10225);
FA fa3286(p10106,p10213,p10092,p10226,p10227);
HA ha1827(p10094,p10096,p10228,p10229);
FA fa3287(p10211,p10215,p10217,p10230,p10231);
HA ha1828(p10219,p10221,p10232,p10233);
HA ha1829(p10223,p10225,p10234,p10235);
FA fa3288(p10100,p10104,p10108,p10236,p10237);
HA ha1830(p10116,p10227,p10238,p10239);
FA fa3289(p10229,p10233,p10235,p10240,p10241);
FA fa3290(p10110,p10112,p10114,p10242,p10243);
HA ha1831(p10231,p10239,p10244,p10245);
FA fa3291(p10118,p10120,p10130,p10246,p10247);
FA fa3292(p10237,p10241,p10245,p10248,p10249);
HA ha1832(p10122,p10124,p10250,p10251);
FA fa3293(p10126,p10128,p10243,p10252,p10253);
HA ha1833(p10132,p10247,p10254,p10255);
FA fa3294(p10249,p10251,p10134,p10256,p10257);
FA fa3295(p10136,p10138,p10142,p10258,p10259);
HA ha1834(p10253,p10255,p10260,p10261);
FA fa3296(p10146,p10257,p10261,p10262,p10263);
HA ha1835(p10140,p10144,p10264,p10265);
FA fa3297(p10259,p10148,p10263,p10266,p10267);
HA ha1836(p10265,p10150,p10268,p10269);
HA ha1837(p10152,p10156,p10270,p10271);
HA ha1838(p10267,p10269,p10272,p10273);
FA fa3298(p10154,p10271,p10273,p10274,p10275);
HA ha1839(p10158,p10275,p10276,p10277);
HA ha1840(p10160,p10277,p10278,p10279);
HA ha1841(p10279,p10162,p10280,p10281);
FA fa3299(ip_30_63,ip_31_62,ip_32_61,p10282,p10283);
HA ha1842(ip_33_60,ip_34_59,p10284,p10285);
FA fa3300(ip_35_58,ip_36_57,ip_37_56,p10286,p10287);
HA ha1843(ip_38_55,ip_39_54,p10288,p10289);
HA ha1844(ip_40_53,ip_41_52,p10290,p10291);
FA fa3301(ip_42_51,ip_43_50,ip_44_49,p10292,p10293);
HA ha1845(ip_45_48,ip_46_47,p10294,p10295);
FA fa3302(ip_47_46,ip_48_45,ip_49_44,p10296,p10297);
FA fa3303(ip_50_43,ip_51_42,ip_52_41,p10298,p10299);
FA fa3304(ip_53_40,ip_54_39,ip_55_38,p10300,p10301);
HA ha1846(ip_56_37,ip_57_36,p10302,p10303);
FA fa3305(ip_58_35,ip_59_34,ip_60_33,p10304,p10305);
FA fa3306(ip_61_32,ip_62_31,ip_63_30,p10306,p10307);
FA fa3307(p10170,p10172,p10178,p10308,p10309);
FA fa3308(p10182,p10184,p10285,p10310,p10311);
FA fa3309(p10289,p10291,p10295,p10312,p10313);
HA ha1847(p10303,p10196,p10314,p10315);
HA ha1848(p10198,p10283,p10316,p10317);
FA fa3310(p10287,p10293,p10297,p10318,p10319);
HA ha1849(p10299,p10301,p10320,p10321);
HA ha1850(p10305,p10307,p10322,p10323);
HA ha1851(p10166,p10168,p10324,p10325);
FA fa3311(p10174,p10176,p10180,p10326,p10327);
FA fa3312(p10186,p10188,p10190,p10328,p10329);
HA ha1852(p10202,p10204,p10330,p10331);
FA fa3313(p10206,p10208,p10309,p10332,p10333);
FA fa3314(p10311,p10313,p10315,p10334,p10335);
FA fa3315(p10317,p10321,p10323,p10336,p10337);
HA ha1853(p10192,p10194,p10338,p10339);
FA fa3316(p10200,p10212,p10319,p10340,p10341);
HA ha1854(p10325,p10331,p10342,p10343);
FA fa3317(p10222,p10224,p10327,p10344,p10345);
FA fa3318(p10329,p10333,p10335,p10346,p10347);
FA fa3319(p10337,p10339,p10343,p10348,p10349);
FA fa3320(p10210,p10214,p10216,p10350,p10351);
HA ha1855(p10218,p10220,p10352,p10353);
FA fa3321(p10228,p10232,p10234,p10354,p10355);
FA fa3322(p10341,p10226,p10238,p10356,p10357);
HA ha1856(p10345,p10347,p10358,p10359);
FA fa3323(p10349,p10353,p10230,p10360,p10361);
FA fa3324(p10244,p10351,p10355,p10362,p10363);
HA ha1857(p10359,p10236,p10364,p10365);
FA fa3325(p10240,p10357,p10361,p10366,p10367);
HA ha1858(p10242,p10250,p10368,p10369);
FA fa3326(p10363,p10365,p10246,p10370,p10371);
HA ha1859(p10248,p10254,p10372,p10373);
FA fa3327(p10367,p10369,p10252,p10374,p10375);
FA fa3328(p10260,p10371,p10373,p10376,p10377);
FA fa3329(p10256,p10375,p10258,p10378,p10379);
FA fa3330(p10264,p10377,p10262,p10380,p10381);
FA fa3331(p10379,p10268,p10381,p10382,p10383);
FA fa3332(p10266,p10270,p10272,p10384,p10385);
FA fa3333(p10383,p10385,p10274,p10386,p10387);
HA ha1860(p10276,p10278,p10388,p10389);
FA fa3334(p10387,p10389,p10280,p10390,p10391);
HA ha1861(ip_31_63,ip_32_62,p10392,p10393);
FA fa3335(ip_33_61,ip_34_60,ip_35_59,p10394,p10395);
FA fa3336(ip_36_58,ip_37_57,ip_38_56,p10396,p10397);
HA ha1862(ip_39_55,ip_40_54,p10398,p10399);
FA fa3337(ip_41_53,ip_42_52,ip_43_51,p10400,p10401);
HA ha1863(ip_44_50,ip_45_49,p10402,p10403);
HA ha1864(ip_46_48,ip_47_47,p10404,p10405);
HA ha1865(ip_48_46,ip_49_45,p10406,p10407);
FA fa3338(ip_50_44,ip_51_43,ip_52_42,p10408,p10409);
FA fa3339(ip_53_41,ip_54_40,ip_55_39,p10410,p10411);
FA fa3340(ip_56_38,ip_57_37,ip_58_36,p10412,p10413);
FA fa3341(ip_59_35,ip_60_34,ip_61_33,p10414,p10415);
FA fa3342(ip_62_32,ip_63_31,p10284,p10416,p10417);
FA fa3343(p10288,p10290,p10294,p10418,p10419);
FA fa3344(p10302,p10393,p10399,p10420,p10421);
HA ha1866(p10403,p10405,p10422,p10423);
FA fa3345(p10407,p10395,p10397,p10424,p10425);
HA ha1867(p10401,p10409,p10426,p10427);
FA fa3346(p10411,p10413,p10415,p10428,p10429);
FA fa3347(p10417,p10423,p10282,p10430,p10431);
HA ha1868(p10286,p10292,p10432,p10433);
FA fa3348(p10296,p10298,p10300,p10434,p10435);
HA ha1869(p10304,p10306,p10436,p10437);
FA fa3349(p10314,p10316,p10320,p10438,p10439);
FA fa3350(p10322,p10419,p10421,p10440,p10441);
FA fa3351(p10427,p10308,p10310,p10442,p10443);
FA fa3352(p10312,p10324,p10330,p10444,p10445);
FA fa3353(p10425,p10429,p10431,p10446,p10447);
FA fa3354(p10433,p10437,p10318,p10448,p10449);
FA fa3355(p10338,p10342,p10435,p10450,p10451);
FA fa3356(p10439,p10441,p10326,p10452,p10453);
FA fa3357(p10328,p10332,p10334,p10454,p10455);
FA fa3358(p10336,p10443,p10445,p10456,p10457);
HA ha1870(p10447,p10449,p10458,p10459);
FA fa3359(p10340,p10352,p10451,p10460,p10461);
HA ha1871(p10453,p10459,p10462,p10463);
FA fa3360(p10344,p10346,p10348,p10464,p10465);
FA fa3361(p10358,p10455,p10457,p10466,p10467);
FA fa3362(p10463,p10350,p10354,p10468,p10469);
FA fa3363(p10461,p10356,p10360,p10470,p10471);
FA fa3364(p10364,p10465,p10467,p10472,p10473);
HA ha1872(p10362,p10368,p10474,p10475);
HA ha1873(p10469,p10366,p10476,p10477);
HA ha1874(p10372,p10471,p10478,p10479);
FA fa3365(p10473,p10475,p10370,p10480,p10481);
FA fa3366(p10477,p10479,p10374,p10482,p10483);
FA fa3367(p10481,p10376,p10483,p10484,p10485);
HA ha1875(p10378,p10380,p10486,p10487);
HA ha1876(p10485,p10487,p10488,p10489);
HA ha1877(p10382,p10489,p10490,p10491);
HA ha1878(p10384,p10491,p10492,p10493);
FA fa3368(p10493,p10386,p10388,p10494,p10495);
HA ha1879(ip_32_63,ip_33_62,p10496,p10497);
HA ha1880(ip_34_61,ip_35_60,p10498,p10499);
FA fa3369(ip_36_59,ip_37_58,ip_38_57,p10500,p10501);
HA ha1881(ip_39_56,ip_40_55,p10502,p10503);
HA ha1882(ip_41_54,ip_42_53,p10504,p10505);
FA fa3370(ip_43_52,ip_44_51,ip_45_50,p10506,p10507);
HA ha1883(ip_46_49,ip_47_48,p10508,p10509);
FA fa3371(ip_48_47,ip_49_46,ip_50_45,p10510,p10511);
FA fa3372(ip_51_44,ip_52_43,ip_53_42,p10512,p10513);
FA fa3373(ip_54_41,ip_55_40,ip_56_39,p10514,p10515);
FA fa3374(ip_57_38,ip_58_37,ip_59_36,p10516,p10517);
HA ha1884(ip_60_35,ip_61_34,p10518,p10519);
HA ha1885(ip_62_33,ip_63_32,p10520,p10521);
FA fa3375(p10392,p10398,p10402,p10522,p10523);
FA fa3376(p10404,p10406,p10497,p10524,p10525);
FA fa3377(p10499,p10503,p10505,p10526,p10527);
HA ha1886(p10509,p10519,p10528,p10529);
FA fa3378(p10521,p10422,p10501,p10530,p10531);
HA ha1887(p10507,p10511,p10532,p10533);
HA ha1888(p10513,p10515,p10534,p10535);
FA fa3379(p10517,p10529,p10394,p10536,p10537);
FA fa3380(p10396,p10400,p10408,p10538,p10539);
FA fa3381(p10410,p10412,p10414,p10540,p10541);
HA ha1889(p10416,p10426,p10542,p10543);
FA fa3382(p10523,p10525,p10527,p10544,p10545);
FA fa3383(p10533,p10535,p10418,p10546,p10547);
HA ha1890(p10420,p10432,p10548,p10549);
HA ha1891(p10436,p10531,p10550,p10551);
HA ha1892(p10537,p10543,p10552,p10553);
FA fa3384(p10424,p10428,p10430,p10554,p10555);
FA fa3385(p10539,p10541,p10545,p10556,p10557);
FA fa3386(p10547,p10549,p10551,p10558,p10559);
HA ha1893(p10553,p10434,p10560,p10561);
HA ha1894(p10438,p10440,p10562,p10563);
FA fa3387(p10442,p10444,p10446,p10564,p10565);
FA fa3388(p10448,p10458,p10555,p10566,p10567);
FA fa3389(p10557,p10559,p10561,p10568,p10569);
HA ha1895(p10563,p10450,p10570,p10571);
HA ha1896(p10452,p10462,p10572,p10573);
HA ha1897(p10454,p10456,p10574,p10575);
FA fa3390(p10565,p10567,p10569,p10576,p10577);
HA ha1898(p10571,p10573,p10578,p10579);
HA ha1899(p10460,p10575,p10580,p10581);
FA fa3391(p10579,p10464,p10466,p10582,p10583);
HA ha1900(p10577,p10581,p10584,p10585);
FA fa3392(p10468,p10474,p10585,p10586,p10587);
FA fa3393(p10470,p10472,p10476,p10588,p10589);
FA fa3394(p10478,p10583,p10587,p10590,p10591);
FA fa3395(p10480,p10589,p10591,p10592,p10593);
FA fa3396(p10482,p10593,p10484,p10594,p10595);
FA fa3397(p10486,p10488,p10595,p10596,p10597);
HA ha1901(p10490,p10492,p10598,p10599);
HA ha1902(p10597,p10599,p10600,p10601);
HA ha1903(ip_33_63,ip_34_62,p10602,p10603);
HA ha1904(ip_35_61,ip_36_60,p10604,p10605);
FA fa3398(ip_37_59,ip_38_58,ip_39_57,p10606,p10607);
HA ha1905(ip_40_56,ip_41_55,p10608,p10609);
HA ha1906(ip_42_54,ip_43_53,p10610,p10611);
FA fa3399(ip_44_52,ip_45_51,ip_46_50,p10612,p10613);
FA fa3400(ip_47_49,ip_48_48,ip_49_47,p10614,p10615);
FA fa3401(ip_50_46,ip_51_45,ip_52_44,p10616,p10617);
FA fa3402(ip_53_43,ip_54_42,ip_55_41,p10618,p10619);
HA ha1907(ip_56_40,ip_57_39,p10620,p10621);
HA ha1908(ip_58_38,ip_59_37,p10622,p10623);
FA fa3403(ip_60_36,ip_61_35,ip_62_34,p10624,p10625);
FA fa3404(ip_63_33,p10496,p10498,p10626,p10627);
FA fa3405(p10502,p10504,p10508,p10628,p10629);
FA fa3406(p10518,p10520,p10603,p10630,p10631);
HA ha1909(p10605,p10609,p10632,p10633);
FA fa3407(p10611,p10621,p10623,p10634,p10635);
HA ha1910(p10528,p10607,p10636,p10637);
HA ha1911(p10613,p10615,p10638,p10639);
HA ha1912(p10617,p10619,p10640,p10641);
FA fa3408(p10625,p10633,p10500,p10642,p10643);
FA fa3409(p10506,p10510,p10512,p10644,p10645);
HA ha1913(p10514,p10516,p10646,p10647);
FA fa3410(p10532,p10534,p10627,p10648,p10649);
HA ha1914(p10629,p10631,p10650,p10651);
FA fa3411(p10635,p10637,p10639,p10652,p10653);
FA fa3412(p10641,p10522,p10524,p10654,p10655);
FA fa3413(p10526,p10542,p10643,p10656,p10657);
FA fa3414(p10647,p10651,p10530,p10658,p10659);
FA fa3415(p10536,p10548,p10550,p10660,p10661);
HA ha1915(p10552,p10645,p10662,p10663);
FA fa3416(p10649,p10653,p10538,p10664,p10665);
FA fa3417(p10540,p10544,p10546,p10666,p10667);
FA fa3418(p10655,p10657,p10659,p10668,p10669);
FA fa3419(p10663,p10560,p10562,p10670,p10671);
FA fa3420(p10661,p10665,p10554,p10672,p10673);
HA ha1916(p10556,p10558,p10674,p10675);
FA fa3421(p10667,p10669,p10570,p10676,p10677);
HA ha1917(p10572,p10671,p10678,p10679);
FA fa3422(p10673,p10675,p10564,p10680,p10681);
HA ha1918(p10566,p10568,p10682,p10683);
FA fa3423(p10574,p10578,p10677,p10684,p10685);
HA ha1919(p10679,p10580,p10686,p10687);
FA fa3424(p10681,p10683,p10576,p10688,p10689);
FA fa3425(p10584,p10685,p10687,p10690,p10691);
FA fa3426(p10689,p10582,p10691,p10692,p10693);
FA fa3427(p10586,p10588,p10590,p10694,p10695);
HA ha1920(p10693,p10592,p10696,p10697);
FA fa3428(p10695,p10697,p10594,p10698,p10699);
FA fa3429(p10699,p10596,p10598,p10700,p10701);
HA ha1921(ip_34_63,ip_35_62,p10702,p10703);
HA ha1922(ip_36_61,ip_37_60,p10704,p10705);
FA fa3430(ip_38_59,ip_39_58,ip_40_57,p10706,p10707);
HA ha1923(ip_41_56,ip_42_55,p10708,p10709);
FA fa3431(ip_43_54,ip_44_53,ip_45_52,p10710,p10711);
HA ha1924(ip_46_51,ip_47_50,p10712,p10713);
FA fa3432(ip_48_49,ip_49_48,ip_50_47,p10714,p10715);
HA ha1925(ip_51_46,ip_52_45,p10716,p10717);
HA ha1926(ip_53_44,ip_54_43,p10718,p10719);
HA ha1927(ip_55_42,ip_56_41,p10720,p10721);
FA fa3433(ip_57_40,ip_58_39,ip_59_38,p10722,p10723);
FA fa3434(ip_60_37,ip_61_36,ip_62_35,p10724,p10725);
HA ha1928(ip_63_34,p10602,p10726,p10727);
FA fa3435(p10604,p10608,p10610,p10728,p10729);
HA ha1929(p10620,p10622,p10730,p10731);
FA fa3436(p10703,p10705,p10709,p10732,p10733);
HA ha1930(p10713,p10717,p10734,p10735);
HA ha1931(p10719,p10721,p10736,p10737);
FA fa3437(p10632,p10707,p10711,p10738,p10739);
FA fa3438(p10715,p10723,p10725,p10740,p10741);
FA fa3439(p10727,p10731,p10735,p10742,p10743);
FA fa3440(p10737,p10606,p10612,p10744,p10745);
HA ha1932(p10614,p10616,p10746,p10747);
FA fa3441(p10618,p10624,p10636,p10748,p10749);
FA fa3442(p10638,p10640,p10729,p10750,p10751);
HA ha1933(p10733,p10626,p10752,p10753);
FA fa3443(p10628,p10630,p10634,p10754,p10755);
FA fa3444(p10646,p10650,p10739,p10756,p10757);
HA ha1934(p10741,p10743,p10758,p10759);
FA fa3445(p10747,p10642,p10745,p10760,p10761);
HA ha1935(p10749,p10751,p10762,p10763);
HA ha1936(p10753,p10759,p10764,p10765);
FA fa3446(p10644,p10648,p10652,p10766,p10767);
FA fa3447(p10662,p10755,p10757,p10768,p10769);
FA fa3448(p10763,p10765,p10654,p10770,p10771);
HA ha1937(p10656,p10658,p10772,p10773);
FA fa3449(p10761,p10660,p10664,p10774,p10775);
HA ha1938(p10767,p10769,p10776,p10777);
FA fa3450(p10771,p10773,p10666,p10778,p10779);
HA ha1939(p10668,p10674,p10780,p10781);
HA ha1940(p10777,p10670,p10782,p10783);
HA ha1941(p10672,p10678,p10784,p10785);
HA ha1942(p10775,p10779,p10786,p10787);
FA fa3451(p10781,p10676,p10682,p10788,p10789);
FA fa3452(p10783,p10785,p10787,p10790,p10791);
FA fa3453(p10680,p10686,p10684,p10792,p10793);
HA ha1943(p10789,p10791,p10794,p10795);
HA ha1944(p10688,p10793,p10796,p10797);
FA fa3454(p10795,p10690,p10797,p10798,p10799);
FA fa3455(p10692,p10799,p10694,p10800,p10801);
HA ha1945(p10696,p10801,p10802,p10803);
HA ha1946(p10803,p10698,p10804,p10805);
FA fa3456(ip_35_63,ip_36_62,ip_37_61,p10806,p10807);
FA fa3457(ip_38_60,ip_39_59,ip_40_58,p10808,p10809);
FA fa3458(ip_41_57,ip_42_56,ip_43_55,p10810,p10811);
FA fa3459(ip_44_54,ip_45_53,ip_46_52,p10812,p10813);
HA ha1947(ip_47_51,ip_48_50,p10814,p10815);
FA fa3460(ip_49_49,ip_50_48,ip_51_47,p10816,p10817);
HA ha1948(ip_52_46,ip_53_45,p10818,p10819);
FA fa3461(ip_54_44,ip_55_43,ip_56_42,p10820,p10821);
FA fa3462(ip_57_41,ip_58_40,ip_59_39,p10822,p10823);
FA fa3463(ip_60_38,ip_61_37,ip_62_36,p10824,p10825);
FA fa3464(ip_63_35,p10702,p10704,p10826,p10827);
FA fa3465(p10708,p10712,p10716,p10828,p10829);
FA fa3466(p10718,p10720,p10815,p10830,p10831);
FA fa3467(p10819,p10726,p10730,p10832,p10833);
FA fa3468(p10734,p10736,p10807,p10834,p10835);
FA fa3469(p10809,p10811,p10813,p10836,p10837);
FA fa3470(p10817,p10821,p10823,p10838,p10839);
FA fa3471(p10825,p10706,p10710,p10840,p10841);
FA fa3472(p10714,p10722,p10724,p10842,p10843);
HA ha1949(p10827,p10829,p10844,p10845);
HA ha1950(p10831,p10728,p10846,p10847);
FA fa3473(p10732,p10746,p10833,p10848,p10849);
FA fa3474(p10835,p10837,p10839,p10850,p10851);
FA fa3475(p10845,p10738,p10740,p10852,p10853);
FA fa3476(p10742,p10752,p10758,p10854,p10855);
FA fa3477(p10841,p10843,p10847,p10856,p10857);
HA ha1951(p10744,p10748,p10858,p10859);
FA fa3478(p10750,p10762,p10764,p10860,p10861);
HA ha1952(p10849,p10851,p10862,p10863);
HA ha1953(p10754,p10756,p10864,p10865);
HA ha1954(p10853,p10855,p10866,p10867);
FA fa3479(p10857,p10859,p10863,p10868,p10869);
HA ha1955(p10760,p10772,p10870,p10871);
FA fa3480(p10861,p10865,p10867,p10872,p10873);
HA ha1956(p10766,p10768,p10874,p10875);
FA fa3481(p10770,p10776,p10869,p10876,p10877);
HA ha1957(p10871,p10780,p10878,p10879);
HA ha1958(p10873,p10875,p10880,p10881);
FA fa3482(p10774,p10778,p10782,p10882,p10883);
HA ha1959(p10784,p10786,p10884,p10885);
HA ha1960(p10877,p10879,p10886,p10887);
HA ha1961(p10881,p10885,p10888,p10889);
FA fa3483(p10887,p10883,p10889,p10890,p10891);
FA fa3484(p10788,p10790,p10794,p10892,p10893);
FA fa3485(p10792,p10796,p10891,p10894,p10895);
HA ha1962(p10893,p10895,p10896,p10897);
FA fa3486(p10798,p10897,p10800,p10898,p10899);
HA ha1963(p10802,p10899,p10900,p10901);
FA fa3487(ip_36_63,ip_37_62,ip_38_61,p10902,p10903);
HA ha1964(ip_39_60,ip_40_59,p10904,p10905);
HA ha1965(ip_41_58,ip_42_57,p10906,p10907);
FA fa3488(ip_43_56,ip_44_55,ip_45_54,p10908,p10909);
HA ha1966(ip_46_53,ip_47_52,p10910,p10911);
FA fa3489(ip_48_51,ip_49_50,ip_50_49,p10912,p10913);
FA fa3490(ip_51_48,ip_52_47,ip_53_46,p10914,p10915);
HA ha1967(ip_54_45,ip_55_44,p10916,p10917);
HA ha1968(ip_56_43,ip_57_42,p10918,p10919);
FA fa3491(ip_58_41,ip_59_40,ip_60_39,p10920,p10921);
HA ha1969(ip_61_38,ip_62_37,p10922,p10923);
FA fa3492(ip_63_36,p10814,p10818,p10924,p10925);
FA fa3493(p10905,p10907,p10911,p10926,p10927);
HA ha1970(p10917,p10919,p10928,p10929);
FA fa3494(p10923,p10903,p10909,p10930,p10931);
HA ha1971(p10913,p10915,p10932,p10933);
FA fa3495(p10921,p10929,p10806,p10934,p10935);
FA fa3496(p10808,p10810,p10812,p10936,p10937);
HA ha1972(p10816,p10820,p10938,p10939);
HA ha1973(p10822,p10824,p10940,p10941);
HA ha1974(p10925,p10927,p10942,p10943);
FA fa3497(p10933,p10826,p10828,p10944,p10945);
HA ha1975(p10830,p10844,p10946,p10947);
FA fa3498(p10931,p10935,p10939,p10948,p10949);
HA ha1976(p10941,p10943,p10950,p10951);
FA fa3499(p10832,p10834,p10836,p10952,p10953);
FA fa3500(p10838,p10846,p10937,p10954,p10955);
FA fa3501(p10947,p10951,p10840,p10956,p10957);
FA fa3502(p10842,p10945,p10949,p10958,p10959);
HA ha1977(p10848,p10850,p10960,p10961);
HA ha1978(p10858,p10862,p10962,p10963);
FA fa3503(p10953,p10955,p10957,p10964,p10965);
FA fa3504(p10852,p10854,p10856,p10966,p10967);
FA fa3505(p10864,p10866,p10959,p10968,p10969);
HA ha1979(p10961,p10963,p10970,p10971);
FA fa3506(p10860,p10870,p10965,p10972,p10973);
FA fa3507(p10971,p10868,p10874,p10974,p10975);
FA fa3508(p10967,p10969,p10872,p10976,p10977);
FA fa3509(p10878,p10880,p10973,p10978,p10979);
FA fa3510(p10876,p10884,p10886,p10980,p10981);
FA fa3511(p10975,p10977,p10888,p10982,p10983);
HA ha1980(p10979,p10882,p10984,p10985);
FA fa3512(p10981,p10983,p10985,p10986,p10987);
FA fa3513(p10890,p10987,p10892,p10988,p10989);
FA fa3514(p10894,p10896,p10989,p10990,p10991);
HA ha1981(p10991,p10898,p10992,p10993);
HA ha1982(ip_37_63,ip_38_62,p10994,p10995);
FA fa3515(ip_39_61,ip_40_60,ip_41_59,p10996,p10997);
FA fa3516(ip_42_58,ip_43_57,ip_44_56,p10998,p10999);
HA ha1983(ip_45_55,ip_46_54,p11000,p11001);
HA ha1984(ip_47_53,ip_48_52,p11002,p11003);
FA fa3517(ip_49_51,ip_50_50,ip_51_49,p11004,p11005);
HA ha1985(ip_52_48,ip_53_47,p11006,p11007);
FA fa3518(ip_54_46,ip_55_45,ip_56_44,p11008,p11009);
FA fa3519(ip_57_43,ip_58_42,ip_59_41,p11010,p11011);
FA fa3520(ip_60_40,ip_61_39,ip_62_38,p11012,p11013);
FA fa3521(ip_63_37,p10904,p10906,p11014,p11015);
HA ha1986(p10910,p10916,p11016,p11017);
FA fa3522(p10918,p10922,p10995,p11018,p11019);
FA fa3523(p11001,p11003,p11007,p11020,p11021);
FA fa3524(p10928,p10997,p10999,p11022,p11023);
HA ha1987(p11005,p11009,p11024,p11025);
FA fa3525(p11011,p11013,p11017,p11026,p11027);
FA fa3526(p10902,p10908,p10912,p11028,p11029);
FA fa3527(p10914,p10920,p10932,p11030,p11031);
FA fa3528(p11015,p11019,p11021,p11032,p11033);
FA fa3529(p11025,p10924,p10926,p11034,p11035);
HA ha1988(p10938,p10940,p11036,p11037);
FA fa3530(p10942,p11023,p11027,p11038,p11039);
FA fa3531(p10930,p10934,p10946,p11040,p11041);
FA fa3532(p10950,p11029,p11031,p11042,p11043);
FA fa3533(p11033,p11037,p10936,p11044,p11045);
FA fa3534(p11035,p11039,p10944,p11046,p11047);
HA ha1989(p10948,p11041,p11048,p11049);
FA fa3535(p11043,p11045,p10952,p11050,p11051);
HA ha1990(p10954,p10956,p11052,p11053);
FA fa3536(p10960,p10962,p11047,p11054,p11055);
FA fa3537(p11049,p10958,p10970,p11056,p11057);
FA fa3538(p11051,p11053,p10964,p11058,p11059);
FA fa3539(p11055,p10966,p10968,p11060,p11061);
FA fa3540(p11057,p11059,p10972,p11062,p11063);
FA fa3541(p10974,p10976,p11061,p11064,p11065);
FA fa3542(p11063,p10978,p10980,p11066,p11067);
HA ha1991(p10982,p10984,p11068,p11069);
HA ha1992(p11065,p11067,p11070,p11071);
HA ha1993(p11069,p10986,p11072,p11073);
FA fa3543(p11071,p11073,p10988,p11074,p11075);
FA fa3544(p11075,p10990,p10992,p11076,p11077);
FA fa3545(ip_38_63,ip_39_62,ip_40_61,p11078,p11079);
FA fa3546(ip_41_60,ip_42_59,ip_43_58,p11080,p11081);
HA ha1994(ip_44_57,ip_45_56,p11082,p11083);
FA fa3547(ip_46_55,ip_47_54,ip_48_53,p11084,p11085);
FA fa3548(ip_49_52,ip_50_51,ip_51_50,p11086,p11087);
FA fa3549(ip_52_49,ip_53_48,ip_54_47,p11088,p11089);
FA fa3550(ip_55_46,ip_56_45,ip_57_44,p11090,p11091);
FA fa3551(ip_58_43,ip_59_42,ip_60_41,p11092,p11093);
HA ha1995(ip_61_40,ip_62_39,p11094,p11095);
FA fa3552(ip_63_38,p10994,p11000,p11096,p11097);
FA fa3553(p11002,p11006,p11083,p11098,p11099);
HA ha1996(p11095,p11016,p11100,p11101);
HA ha1997(p11079,p11081,p11102,p11103);
FA fa3554(p11085,p11087,p11089,p11104,p11105);
HA ha1998(p11091,p11093,p11106,p11107);
HA ha1999(p10996,p10998,p11108,p11109);
HA ha2000(p11004,p11008,p11110,p11111);
HA ha2001(p11010,p11012,p11112,p11113);
HA ha2002(p11024,p11097,p11114,p11115);
FA fa3555(p11099,p11101,p11103,p11116,p11117);
FA fa3556(p11107,p11014,p11018,p11118,p11119);
FA fa3557(p11020,p11105,p11109,p11120,p11121);
HA ha2003(p11111,p11113,p11122,p11123);
HA ha2004(p11115,p11022,p11124,p11125);
FA fa3558(p11026,p11036,p11117,p11126,p11127);
FA fa3559(p11123,p11028,p11030,p11128,p11129);
FA fa3560(p11032,p11119,p11121,p11130,p11131);
FA fa3561(p11125,p11034,p11038,p11132,p11133);
FA fa3562(p11127,p11040,p11042,p11134,p11135);
FA fa3563(p11044,p11048,p11129,p11136,p11137);
HA ha2005(p11131,p11046,p11138,p11139);
FA fa3564(p11052,p11133,p11050,p11140,p11141);
HA ha2006(p11135,p11137,p11142,p11143);
FA fa3565(p11139,p11054,p11141,p11144,p11145);
FA fa3566(p11143,p11056,p11058,p11146,p11147);
FA fa3567(p11145,p11060,p11062,p11148,p11149);
HA ha2007(p11147,p11064,p11150,p11151);
FA fa3568(p11068,p11149,p11066,p11152,p11153);
FA fa3569(p11070,p11151,p11072,p11154,p11155);
FA fa3570(p11153,p11155,p11074,p11156,p11157);
HA ha2008(ip_39_63,ip_40_62,p11158,p11159);
FA fa3571(ip_41_61,ip_42_60,ip_43_59,p11160,p11161);
FA fa3572(ip_44_58,ip_45_57,ip_46_56,p11162,p11163);
FA fa3573(ip_47_55,ip_48_54,ip_49_53,p11164,p11165);
FA fa3574(ip_50_52,ip_51_51,ip_52_50,p11166,p11167);
HA ha2009(ip_53_49,ip_54_48,p11168,p11169);
HA ha2010(ip_55_47,ip_56_46,p11170,p11171);
FA fa3575(ip_57_45,ip_58_44,ip_59_43,p11172,p11173);
FA fa3576(ip_60_42,ip_61_41,ip_62_40,p11174,p11175);
FA fa3577(ip_63_39,p11082,p11094,p11176,p11177);
HA ha2011(p11159,p11169,p11178,p11179);
HA ha2012(p11171,p11161,p11180,p11181);
FA fa3578(p11163,p11165,p11167,p11182,p11183);
HA ha2013(p11173,p11175,p11184,p11185);
FA fa3579(p11179,p11078,p11080,p11186,p11187);
HA ha2014(p11084,p11086,p11188,p11189);
FA fa3580(p11088,p11090,p11092,p11190,p11191);
FA fa3581(p11100,p11102,p11106,p11192,p11193);
HA ha2015(p11177,p11181,p11194,p11195);
FA fa3582(p11185,p11096,p11098,p11196,p11197);
FA fa3583(p11108,p11110,p11112,p11198,p11199);
HA ha2016(p11114,p11183,p11200,p11201);
HA ha2017(p11189,p11195,p11202,p11203);
FA fa3584(p11104,p11122,p11187,p11204,p11205);
HA ha2018(p11191,p11193,p11206,p11207);
FA fa3585(p11201,p11203,p11116,p11208,p11209);
HA ha2019(p11124,p11197,p11210,p11211);
FA fa3586(p11199,p11207,p11118,p11212,p11213);
HA ha2020(p11120,p11205,p11214,p11215);
FA fa3587(p11209,p11211,p11126,p11216,p11217);
FA fa3588(p11213,p11215,p11128,p11218,p11219);
HA ha2021(p11130,p11217,p11220,p11221);
FA fa3589(p11132,p11138,p11219,p11222,p11223);
FA fa3590(p11221,p11134,p11136,p11224,p11225);
HA ha2022(p11142,p11140,p11226,p11227);
HA ha2023(p11223,p11225,p11228,p11229);
HA ha2024(p11227,p11144,p11230,p11231);
HA ha2025(p11229,p11146,p11232,p11233);
FA fa3591(p11231,p11233,p11148,p11234,p11235);
FA fa3592(p11150,p11235,p11152,p11236,p11237);
FA fa3593(p11154,p11237,p11156,p11238,p11239);
FA fa3594(ip_40_63,ip_41_62,ip_42_61,p11240,p11241);
FA fa3595(ip_43_60,ip_44_59,ip_45_58,p11242,p11243);
FA fa3596(ip_46_57,ip_47_56,ip_48_55,p11244,p11245);
HA ha2026(ip_49_54,ip_50_53,p11246,p11247);
HA ha2027(ip_51_52,ip_52_51,p11248,p11249);
HA ha2028(ip_53_50,ip_54_49,p11250,p11251);
FA fa3597(ip_55_48,ip_56_47,ip_57_46,p11252,p11253);
HA ha2029(ip_58_45,ip_59_44,p11254,p11255);
FA fa3598(ip_60_43,ip_61_42,ip_62_41,p11256,p11257);
FA fa3599(ip_63_40,p11158,p11168,p11258,p11259);
HA ha2030(p11170,p11247,p11260,p11261);
FA fa3600(p11249,p11251,p11255,p11262,p11263);
FA fa3601(p11178,p11241,p11243,p11264,p11265);
FA fa3602(p11245,p11253,p11257,p11266,p11267);
HA ha2031(p11261,p11160,p11268,p11269);
FA fa3603(p11162,p11164,p11166,p11270,p11271);
FA fa3604(p11172,p11174,p11180,p11272,p11273);
HA ha2032(p11184,p11259,p11274,p11275);
HA ha2033(p11263,p11176,p11276,p11277);
FA fa3605(p11188,p11194,p11265,p11278,p11279);
FA fa3606(p11267,p11269,p11275,p11280,p11281);
HA ha2034(p11182,p11200,p11282,p11283);
HA ha2035(p11202,p11271,p11284,p11285);
HA ha2036(p11273,p11277,p11286,p11287);
HA ha2037(p11186,p11190,p11288,p11289);
HA ha2038(p11192,p11206,p11290,p11291);
FA fa3607(p11279,p11281,p11283,p11292,p11293);
FA fa3608(p11285,p11287,p11196,p11294,p11295);
FA fa3609(p11198,p11210,p11289,p11296,p11297);
FA fa3610(p11291,p11204,p11208,p11298,p11299);
FA fa3611(p11214,p11293,p11295,p11300,p11301);
FA fa3612(p11212,p11297,p11216,p11302,p11303);
FA fa3613(p11220,p11299,p11301,p11304,p11305);
FA fa3614(p11218,p11303,p11305,p11306,p11307);
HA ha2039(p11222,p11226,p11308,p11309);
FA fa3615(p11307,p11224,p11228,p11310,p11311);
HA ha2040(p11309,p11230,p11312,p11313);
HA ha2041(p11232,p11311,p11314,p11315);
HA ha2042(p11313,p11315,p11316,p11317);
FA fa3616(p11317,p11234,p11236,p11318,p11319);
FA fa3617(ip_41_63,ip_42_62,ip_43_61,p11320,p11321);
FA fa3618(ip_44_60,ip_45_59,ip_46_58,p11322,p11323);
HA ha2043(ip_47_57,ip_48_56,p11324,p11325);
FA fa3619(ip_49_55,ip_50_54,ip_51_53,p11326,p11327);
HA ha2044(ip_52_52,ip_53_51,p11328,p11329);
HA ha2045(ip_54_50,ip_55_49,p11330,p11331);
FA fa3620(ip_56_48,ip_57_47,ip_58_46,p11332,p11333);
FA fa3621(ip_59_45,ip_60_44,ip_61_43,p11334,p11335);
HA ha2046(ip_62_42,ip_63_41,p11336,p11337);
FA fa3622(p11246,p11248,p11250,p11338,p11339);
HA ha2047(p11254,p11325,p11340,p11341);
FA fa3623(p11329,p11331,p11337,p11342,p11343);
FA fa3624(p11260,p11321,p11323,p11344,p11345);
FA fa3625(p11327,p11333,p11335,p11346,p11347);
FA fa3626(p11341,p11240,p11242,p11348,p11349);
FA fa3627(p11244,p11252,p11256,p11350,p11351);
FA fa3628(p11339,p11343,p11258,p11352,p11353);
FA fa3629(p11262,p11268,p11274,p11354,p11355);
FA fa3630(p11345,p11347,p11264,p11356,p11357);
FA fa3631(p11266,p11276,p11349,p11358,p11359);
FA fa3632(p11351,p11353,p11270,p11360,p11361);
HA ha2048(p11272,p11282,p11362,p11363);
FA fa3633(p11284,p11286,p11355,p11364,p11365);
FA fa3634(p11357,p11278,p11280,p11366,p11367);
FA fa3635(p11288,p11290,p11359,p11368,p11369);
HA ha2049(p11361,p11363,p11370,p11371);
FA fa3636(p11365,p11371,p11292,p11372,p11373);
FA fa3637(p11294,p11367,p11369,p11374,p11375);
FA fa3638(p11296,p11373,p11298,p11376,p11377);
FA fa3639(p11300,p11375,p11302,p11378,p11379);
HA ha2050(p11377,p11304,p11380,p11381);
FA fa3640(p11379,p11306,p11308,p11382,p11383);
HA ha2051(p11381,p11312,p11384,p11385);
FA fa3641(p11383,p11310,p11314,p11386,p11387);
FA fa3642(p11385,p11316,p11387,p11388,p11389);
FA fa3643(ip_42_63,ip_43_62,ip_44_61,p11390,p11391);
HA ha2052(ip_45_60,ip_46_59,p11392,p11393);
FA fa3644(ip_47_58,ip_48_57,ip_49_56,p11394,p11395);
FA fa3645(ip_50_55,ip_51_54,ip_52_53,p11396,p11397);
FA fa3646(ip_53_52,ip_54_51,ip_55_50,p11398,p11399);
HA ha2053(ip_56_49,ip_57_48,p11400,p11401);
FA fa3647(ip_58_47,ip_59_46,ip_60_45,p11402,p11403);
FA fa3648(ip_61_44,ip_62_43,ip_63_42,p11404,p11405);
HA ha2054(p11324,p11328,p11406,p11407);
FA fa3649(p11330,p11336,p11393,p11408,p11409);
HA ha2055(p11401,p11340,p11410,p11411);
HA ha2056(p11391,p11395,p11412,p11413);
FA fa3650(p11397,p11399,p11403,p11414,p11415);
FA fa3651(p11405,p11407,p11320,p11416,p11417);
HA ha2057(p11322,p11326,p11418,p11419);
HA ha2058(p11332,p11334,p11420,p11421);
HA ha2059(p11409,p11411,p11422,p11423);
FA fa3652(p11413,p11338,p11342,p11424,p11425);
FA fa3653(p11415,p11417,p11419,p11426,p11427);
FA fa3654(p11421,p11423,p11344,p11428,p11429);
FA fa3655(p11346,p11348,p11350,p11430,p11431);
FA fa3656(p11352,p11425,p11427,p11432,p11433);
FA fa3657(p11429,p11354,p11356,p11434,p11435);
FA fa3658(p11362,p11358,p11360,p11436,p11437);
FA fa3659(p11370,p11431,p11433,p11438,p11439);
HA ha2060(p11364,p11435,p11440,p11441);
FA fa3660(p11366,p11368,p11437,p11442,p11443);
HA ha2061(p11439,p11441,p11444,p11445);
HA ha2062(p11372,p11445,p11446,p11447);
HA ha2063(p11374,p11443,p11448,p11449);
FA fa3661(p11447,p11376,p11449,p11450,p11451);
FA fa3662(p11378,p11380,p11451,p11452,p11453);
FA fa3663(p11453,p11382,p11384,p11454,p11455);
HA ha2064(p11455,p11386,p11456,p11457);
FA fa3664(ip_43_63,ip_44_62,ip_45_61,p11458,p11459);
FA fa3665(ip_46_60,ip_47_59,ip_48_58,p11460,p11461);
FA fa3666(ip_49_57,ip_50_56,ip_51_55,p11462,p11463);
FA fa3667(ip_52_54,ip_53_53,ip_54_52,p11464,p11465);
FA fa3668(ip_55_51,ip_56_50,ip_57_49,p11466,p11467);
HA ha2065(ip_58_48,ip_59_47,p11468,p11469);
HA ha2066(ip_60_46,ip_61_45,p11470,p11471);
FA fa3669(ip_62_44,ip_63_43,p11392,p11472,p11473);
HA ha2067(p11400,p11469,p11474,p11475);
FA fa3670(p11471,p11406,p11459,p11476,p11477);
HA ha2068(p11461,p11463,p11478,p11479);
FA fa3671(p11465,p11467,p11473,p11480,p11481);
FA fa3672(p11475,p11390,p11394,p11482,p11483);
HA ha2069(p11396,p11398,p11484,p11485);
FA fa3673(p11402,p11404,p11410,p11486,p11487);
FA fa3674(p11412,p11479,p11408,p11488,p11489);
HA ha2070(p11418,p11420,p11490,p11491);
FA fa3675(p11422,p11477,p11481,p11492,p11493);
HA ha2071(p11485,p11414,p11494,p11495);
FA fa3676(p11416,p11483,p11487,p11496,p11497);
FA fa3677(p11489,p11491,p11493,p11498,p11499);
FA fa3678(p11495,p11424,p11426,p11500,p11501);
FA fa3679(p11428,p11497,p11499,p11502,p11503);
FA fa3680(p11430,p11432,p11501,p11504,p11505);
FA fa3681(p11503,p11434,p11440,p11506,p11507);
HA ha2072(p11436,p11438,p11508,p11509);
HA ha2073(p11444,p11505,p11510,p11511);
FA fa3682(p11446,p11507,p11509,p11512,p11513);
HA ha2074(p11511,p11442,p11514,p11515);
HA ha2075(p11448,p11513,p11516,p11517);
FA fa3683(p11515,p11517,p11450,p11518,p11519);
FA fa3684(p11452,p11519,p11454,p11520,p11521);
HA ha2076(ip_44_63,ip_45_62,p11522,p11523);
FA fa3685(ip_46_61,ip_47_60,ip_48_59,p11524,p11525);
FA fa3686(ip_49_58,ip_50_57,ip_51_56,p11526,p11527);
FA fa3687(ip_52_55,ip_53_54,ip_54_53,p11528,p11529);
HA ha2077(ip_55_52,ip_56_51,p11530,p11531);
HA ha2078(ip_57_50,ip_58_49,p11532,p11533);
HA ha2079(ip_59_48,ip_60_47,p11534,p11535);
HA ha2080(ip_61_46,ip_62_45,p11536,p11537);
FA fa3688(ip_63_44,p11468,p11470,p11538,p11539);
HA ha2081(p11523,p11531,p11540,p11541);
HA ha2082(p11533,p11535,p11542,p11543);
HA ha2083(p11537,p11474,p11544,p11545);
HA ha2084(p11525,p11527,p11546,p11547);
FA fa3689(p11529,p11541,p11543,p11548,p11549);
HA ha2085(p11458,p11460,p11550,p11551);
FA fa3690(p11462,p11464,p11466,p11552,p11553);
FA fa3691(p11472,p11478,p11539,p11554,p11555);
HA ha2086(p11545,p11547,p11556,p11557);
FA fa3692(p11484,p11549,p11551,p11558,p11559);
FA fa3693(p11557,p11476,p11480,p11560,p11561);
FA fa3694(p11490,p11553,p11555,p11562,p11563);
HA ha2087(p11482,p11486,p11564,p11565);
FA fa3695(p11488,p11494,p11559,p11566,p11567);
FA fa3696(p11492,p11561,p11563,p11568,p11569);
FA fa3697(p11565,p11496,p11498,p11570,p11571);
HA ha2088(p11567,p11569,p11572,p11573);
FA fa3698(p11500,p11502,p11571,p11574,p11575);
FA fa3699(p11573,p11504,p11508,p11576,p11577);
FA fa3700(p11510,p11575,p11506,p11578,p11579);
FA fa3701(p11514,p11577,p11579,p11580,p11581);
HA ha2089(p11512,p11516,p11582,p11583);
HA ha2090(p11581,p11583,p11584,p11585);
FA fa3702(p11585,p11518,p11520,p11586,p11587);
HA ha2091(ip_45_63,ip_46_62,p11588,p11589);
HA ha2092(ip_47_61,ip_48_60,p11590,p11591);
FA fa3703(ip_49_59,ip_50_58,ip_51_57,p11592,p11593);
FA fa3704(ip_52_56,ip_53_55,ip_54_54,p11594,p11595);
FA fa3705(ip_55_53,ip_56_52,ip_57_51,p11596,p11597);
HA ha2093(ip_58_50,ip_59_49,p11598,p11599);
HA ha2094(ip_60_48,ip_61_47,p11600,p11601);
HA ha2095(ip_62_46,ip_63_45,p11602,p11603);
HA ha2096(p11522,p11530,p11604,p11605);
FA fa3706(p11532,p11534,p11536,p11606,p11607);
FA fa3707(p11589,p11591,p11599,p11608,p11609);
HA ha2097(p11601,p11603,p11610,p11611);
FA fa3708(p11540,p11542,p11593,p11612,p11613);
FA fa3709(p11595,p11597,p11605,p11614,p11615);
FA fa3710(p11611,p11524,p11526,p11616,p11617);
HA ha2098(p11528,p11544,p11618,p11619);
FA fa3711(p11546,p11607,p11609,p11620,p11621);
HA ha2099(p11538,p11550,p11622,p11623);
FA fa3712(p11556,p11613,p11615,p11624,p11625);
FA fa3713(p11619,p11548,p11617,p11626,p11627);
FA fa3714(p11621,p11623,p11552,p11628,p11629);
HA ha2100(p11554,p11625,p11630,p11631);
FA fa3715(p11558,p11564,p11627,p11632,p11633);
FA fa3716(p11629,p11631,p11560,p11634,p11635);
FA fa3717(p11562,p11566,p11633,p11636,p11637);
FA fa3718(p11635,p11568,p11572,p11638,p11639);
FA fa3719(p11570,p11637,p11639,p11640,p11641);
FA fa3720(p11574,p11641,p11576,p11642,p11643);
FA fa3721(p11578,p11582,p11643,p11644,p11645);
HA ha2101(p11580,p11584,p11646,p11647);
FA fa3722(p11645,p11647,p11586,p11648,p11649);
HA ha2102(ip_46_63,ip_47_62,p11650,p11651);
FA fa3723(ip_48_61,ip_49_60,ip_50_59,p11652,p11653);
FA fa3724(ip_51_58,ip_52_57,ip_53_56,p11654,p11655);
FA fa3725(ip_54_55,ip_55_54,ip_56_53,p11656,p11657);
FA fa3726(ip_57_52,ip_58_51,ip_59_50,p11658,p11659);
FA fa3727(ip_60_49,ip_61_48,ip_62_47,p11660,p11661);
FA fa3728(ip_63_46,p11588,p11590,p11662,p11663);
FA fa3729(p11598,p11600,p11602,p11664,p11665);
HA ha2103(p11651,p11604,p11666,p11667);
HA ha2104(p11610,p11653,p11668,p11669);
HA ha2105(p11655,p11657,p11670,p11671);
HA ha2106(p11659,p11661,p11672,p11673);
HA ha2107(p11592,p11594,p11674,p11675);
FA fa3730(p11596,p11663,p11665,p11676,p11677);
HA ha2108(p11667,p11669,p11678,p11679);
FA fa3731(p11671,p11673,p11606,p11680,p11681);
FA fa3732(p11608,p11618,p11675,p11682,p11683);
FA fa3733(p11679,p11612,p11614,p11684,p11685);
FA fa3734(p11622,p11677,p11681,p11686,p11687);
FA fa3735(p11616,p11620,p11683,p11688,p11689);
FA fa3736(p11624,p11630,p11685,p11690,p11691);
FA fa3737(p11687,p11626,p11628,p11692,p11693);
FA fa3738(p11689,p11691,p11632,p11694,p11695);
FA fa3739(p11634,p11693,p11695,p11696,p11697);
FA fa3740(p11636,p11697,p11638,p11698,p11699);
FA fa3741(p11640,p11699,p11642,p11700,p11701);
FA fa3742(p11646,p11701,p11644,p11702,p11703);
FA fa3743(ip_47_63,ip_48_62,ip_49_61,p11704,p11705);
FA fa3744(ip_50_60,ip_51_59,ip_52_58,p11706,p11707);
HA ha2109(ip_53_57,ip_54_56,p11708,p11709);
HA ha2110(ip_55_55,ip_56_54,p11710,p11711);
HA ha2111(ip_57_53,ip_58_52,p11712,p11713);
FA fa3745(ip_59_51,ip_60_50,ip_61_49,p11714,p11715);
HA ha2112(ip_62_48,ip_63_47,p11716,p11717);
HA ha2113(p11650,p11709,p11718,p11719);
FA fa3746(p11711,p11713,p11717,p11720,p11721);
HA ha2114(p11705,p11707,p11722,p11723);
FA fa3747(p11715,p11719,p11652,p11724,p11725);
HA ha2115(p11654,p11656,p11726,p11727);
FA fa3748(p11658,p11660,p11666,p11728,p11729);
FA fa3749(p11668,p11670,p11672,p11730,p11731);
HA ha2116(p11721,p11723,p11732,p11733);
HA ha2117(p11662,p11664,p11734,p11735);
HA ha2118(p11674,p11678,p11736,p11737);
HA ha2119(p11725,p11727,p11738,p11739);
HA ha2120(p11733,p11729,p11740,p11741);
HA ha2121(p11731,p11735,p11742,p11743);
FA fa3750(p11737,p11739,p11676,p11744,p11745);
FA fa3751(p11680,p11741,p11743,p11746,p11747);
FA fa3752(p11682,p11745,p11684,p11748,p11749);
HA ha2122(p11686,p11747,p11750,p11751);
FA fa3753(p11688,p11749,p11751,p11752,p11753);
FA fa3754(p11690,p11692,p11753,p11754,p11755);
HA ha2123(p11694,p11696,p11756,p11757);
HA ha2124(p11755,p11757,p11758,p11759);
HA ha2125(p11698,p11759,p11760,p11761);
FA fa3755(p11761,p11700,p11702,p11762,p11763);
FA fa3756(ip_48_63,ip_49_62,ip_50_61,p11764,p11765);
FA fa3757(ip_51_60,ip_52_59,ip_53_58,p11766,p11767);
HA ha2126(ip_54_57,ip_55_56,p11768,p11769);
HA ha2127(ip_56_55,ip_57_54,p11770,p11771);
HA ha2128(ip_58_53,ip_59_52,p11772,p11773);
FA fa3758(ip_60_51,ip_61_50,ip_62_49,p11774,p11775);
HA ha2129(ip_63_48,p11708,p11776,p11777);
FA fa3759(p11710,p11712,p11716,p11778,p11779);
FA fa3760(p11769,p11771,p11773,p11780,p11781);
FA fa3761(p11718,p11765,p11767,p11782,p11783);
FA fa3762(p11775,p11777,p11704,p11784,p11785);
FA fa3763(p11706,p11714,p11722,p11786,p11787);
HA ha2130(p11779,p11781,p11788,p11789);
FA fa3764(p11720,p11726,p11732,p11790,p11791);
FA fa3765(p11783,p11785,p11789,p11792,p11793);
FA fa3766(p11724,p11734,p11736,p11794,p11795);
FA fa3767(p11738,p11787,p11728,p11796,p11797);
HA ha2131(p11730,p11740,p11798,p11799);
FA fa3768(p11742,p11791,p11793,p11800,p11801);
FA fa3769(p11795,p11797,p11799,p11802,p11803);
FA fa3770(p11744,p11801,p11746,p11804,p11805);
FA fa3771(p11750,p11803,p11748,p11806,p11807);
FA fa3772(p11805,p11807,p11752,p11808,p11809);
HA ha2132(p11809,p11754,p11810,p11811);
HA ha2133(p11756,p11758,p11812,p11813);
FA fa3773(p11811,p11760,p11813,p11814,p11815);
HA ha2134(ip_49_63,ip_50_62,p11816,p11817);
FA fa3774(ip_51_61,ip_52_60,ip_53_59,p11818,p11819);
HA ha2135(ip_54_58,ip_55_57,p11820,p11821);
HA ha2136(ip_56_56,ip_57_55,p11822,p11823);
HA ha2137(ip_58_54,ip_59_53,p11824,p11825);
FA fa3775(ip_60_52,ip_61_51,ip_62_50,p11826,p11827);
FA fa3776(ip_63_49,p11768,p11770,p11828,p11829);
FA fa3777(p11772,p11817,p11821,p11830,p11831);
FA fa3778(p11823,p11825,p11776,p11832,p11833);
HA ha2138(p11819,p11827,p11834,p11835);
FA fa3779(p11764,p11766,p11774,p11836,p11837);
FA fa3780(p11829,p11831,p11833,p11838,p11839);
FA fa3781(p11835,p11778,p11780,p11840,p11841);
FA fa3782(p11788,p11782,p11784,p11842,p11843);
FA fa3783(p11837,p11839,p11786,p11844,p11845);
FA fa3784(p11841,p11790,p11792,p11846,p11847);
HA ha2139(p11798,p11843,p11848,p11849);
FA fa3785(p11845,p11794,p11796,p11850,p11851);
FA fa3786(p11849,p11800,p11847,p11852,p11853);
HA ha2140(p11802,p11851,p11854,p11855);
FA fa3787(p11804,p11853,p11855,p11856,p11857);
FA fa3788(p11806,p11857,p11808,p11858,p11859);
FA fa3789(p11810,p11859,p11812,p11860,p11861);
FA fa3790(ip_50_63,ip_51_62,ip_52_61,p11862,p11863);
HA ha2141(ip_53_60,ip_54_59,p11864,p11865);
FA fa3791(ip_55_58,ip_56_57,ip_57_56,p11866,p11867);
FA fa3792(ip_58_55,ip_59_54,ip_60_53,p11868,p11869);
FA fa3793(ip_61_52,ip_62_51,ip_63_50,p11870,p11871);
HA ha2142(p11816,p11820,p11872,p11873);
HA ha2143(p11822,p11824,p11874,p11875);
HA ha2144(p11865,p11863,p11876,p11877);
FA fa3794(p11867,p11869,p11871,p11878,p11879);
FA fa3795(p11873,p11875,p11818,p11880,p11881);
FA fa3796(p11826,p11834,p11877,p11882,p11883);
FA fa3797(p11828,p11830,p11832,p11884,p11885);
FA fa3798(p11879,p11881,p11883,p11886,p11887);
FA fa3799(p11836,p11838,p11885,p11888,p11889);
HA ha2145(p11887,p11840,p11890,p11891);
FA fa3800(p11842,p11844,p11848,p11892,p11893);
FA fa3801(p11889,p11891,p11846,p11894,p11895);
FA fa3802(p11893,p11850,p11854,p11896,p11897);
HA ha2146(p11895,p11852,p11898,p11899);
FA fa3803(p11897,p11899,p11856,p11900,p11901);
HA ha2147(p11901,p11858,p11902,p11903);
FA fa3804(ip_51_63,ip_52_62,ip_53_61,p11904,p11905);
FA fa3805(ip_54_60,ip_55_59,ip_56_58,p11906,p11907);
FA fa3806(ip_57_57,ip_58_56,ip_59_55,p11908,p11909);
FA fa3807(ip_60_54,ip_61_53,ip_62_52,p11910,p11911);
FA fa3808(ip_63_51,p11864,p11872,p11912,p11913);
HA ha2148(p11874,p11905,p11914,p11915);
HA ha2149(p11907,p11909,p11916,p11917);
FA fa3809(p11911,p11862,p11866,p11918,p11919);
FA fa3810(p11868,p11870,p11876,p11920,p11921);
FA fa3811(p11913,p11915,p11917,p11922,p11923);
FA fa3812(p11878,p11880,p11919,p11924,p11925);
HA ha2150(p11921,p11923,p11926,p11927);
HA ha2151(p11882,p11927,p11928,p11929);
FA fa3813(p11884,p11886,p11925,p11930,p11931);
FA fa3814(p11929,p11890,p11888,p11932,p11933);
FA fa3815(p11931,p11933,p11892,p11934,p11935);
FA fa3816(p11894,p11935,p11898,p11936,p11937);
FA fa3817(p11896,p11937,p11900,p11938,p11939);
HA ha2152(ip_52_63,ip_53_62,p11940,p11941);
FA fa3818(ip_54_61,ip_55_60,ip_56_59,p11942,p11943);
FA fa3819(ip_57_58,ip_58_57,ip_59_56,p11944,p11945);
FA fa3820(ip_60_55,ip_61_54,ip_62_53,p11946,p11947);
FA fa3821(ip_63_52,p11941,p11943,p11948,p11949);
FA fa3822(p11945,p11947,p11904,p11950,p11951);
FA fa3823(p11906,p11908,p11910,p11952,p11953);
HA ha2153(p11914,p11916,p11954,p11955);
FA fa3824(p11949,p11912,p11951,p11956,p11957);
FA fa3825(p11955,p11953,p11918,p11958,p11959);
HA ha2154(p11920,p11922,p11960,p11961);
FA fa3826(p11926,p11957,p11928,p11962,p11963);
HA ha2155(p11959,p11961,p11964,p11965);
HA ha2156(p11924,p11963,p11966,p11967);
FA fa3827(p11965,p11967,p11930,p11968,p11969);
FA fa3828(p11932,p11969,p11934,p11970,p11971);
FA fa3829(p11971,p11936,p11938,p11972,p11973);
FA fa3830(ip_53_63,ip_54_62,ip_55_61,p11974,p11975);
HA ha2157(ip_56_60,ip_57_59,p11976,p11977);
FA fa3831(ip_58_58,ip_59_57,ip_60_56,p11978,p11979);
FA fa3832(ip_61_55,ip_62_54,ip_63_53,p11980,p11981);
FA fa3833(p11940,p11977,p11975,p11982,p11983);
HA ha2158(p11979,p11981,p11984,p11985);
FA fa3834(p11942,p11944,p11946,p11986,p11987);
FA fa3835(p11983,p11985,p11948,p11988,p11989);
FA fa3836(p11954,p11950,p11987,p11990,p11991);
FA fa3837(p11989,p11952,p11956,p11992,p11993);
FA fa3838(p11960,p11991,p11958,p11994,p11995);
HA ha2159(p11964,p11993,p11996,p11997);
FA fa3839(p11962,p11966,p11995,p11998,p11999);
FA fa3840(p11997,p11999,p11968,p12000,p12001);
HA ha2160(p12001,p11970,p12002,p12003);
FA fa3841(ip_54_63,ip_55_62,ip_56_61,p12004,p12005);
HA ha2161(ip_57_60,ip_58_59,p12006,p12007);
HA ha2162(ip_59_58,ip_60_57,p12008,p12009);
FA fa3842(ip_61_56,ip_62_55,ip_63_54,p12010,p12011);
HA ha2163(p11976,p12007,p12012,p12013);
FA fa3843(p12009,p12005,p12011,p12014,p12015);
HA ha2164(p12013,p11974,p12016,p12017);
HA ha2165(p11978,p11980,p12018,p12019);
FA fa3844(p11984,p11982,p12015,p12020,p12021);
FA fa3845(p12017,p12019,p11986,p12022,p12023);
HA ha2166(p11988,p12021,p12024,p12025);
FA fa3846(p12023,p12025,p11990,p12026,p12027);
HA ha2167(p11992,p11996,p12028,p12029);
FA fa3847(p12027,p11994,p12029,p12030,p12031);
FA fa3848(p11998,p12031,p12000,p12032,p12033);
HA ha2168(ip_55_63,ip_56_62,p12034,p12035);
FA fa3849(ip_57_61,ip_58_60,ip_59_59,p12036,p12037);
HA ha2169(ip_60_58,ip_61_57,p12038,p12039);
HA ha2170(ip_62_56,ip_63_55,p12040,p12041);
FA fa3850(p12006,p12008,p12035,p12042,p12043);
HA ha2171(p12039,p12041,p12044,p12045);
HA ha2172(p12012,p12037,p12046,p12047);
HA ha2173(p12045,p12004,p12048,p12049);
FA fa3851(p12010,p12043,p12047,p12050,p12051);
FA fa3852(p12016,p12018,p12049,p12052,p12053);
FA fa3853(p12014,p12051,p12053,p12054,p12055);
FA fa3854(p12020,p12024,p12055,p12056,p12057);
FA fa3855(p12022,p12057,p12026,p12058,p12059);
FA fa3856(p12028,p12059,p12030,p12060,p12061);
FA fa3857(ip_56_63,ip_57_62,ip_58_61,p12062,p12063);
FA fa3858(ip_59_60,ip_60_59,ip_61_58,p12064,p12065);
HA ha2174(ip_62_57,ip_63_56,p12066,p12067);
FA fa3859(p12034,p12038,p12040,p12068,p12069);
FA fa3860(p12067,p12044,p12063,p12070,p12071);
FA fa3861(p12065,p12036,p12046,p12072,p12073);
HA ha2175(p12069,p12042,p12074,p12075);
HA ha2176(p12048,p12071,p12076,p12077);
HA ha2177(p12073,p12075,p12078,p12079);
HA ha2178(p12077,p12050,p12080,p12081);
FA fa3862(p12079,p12052,p12081,p12082,p12083);
FA fa3863(p12054,p12083,p12056,p12084,p12085);
HA ha2179(p12085,p12058,p12086,p12087);
FA fa3864(ip_57_63,ip_58_62,ip_59_61,p12088,p12089);
FA fa3865(ip_60_60,ip_61_59,ip_62_58,p12090,p12091);
HA ha2180(ip_63_57,p12066,p12092,p12093);
HA ha2181(p12089,p12091,p12094,p12095);
HA ha2182(p12093,p12062,p12096,p12097);
HA ha2183(p12064,p12095,p12098,p12099);
HA ha2184(p12068,p12097,p12100,p12101);
FA fa3866(p12099,p12070,p12074,p12102,p12103);
FA fa3867(p12076,p12101,p12072,p12104,p12105);
HA ha2185(p12078,p12080,p12106,p12107);
FA fa3868(p12103,p12105,p12107,p12108,p12109);
FA fa3869(p12109,p12082,p12084,p12110,p12111);
HA ha2186(ip_58_63,ip_59_62,p12112,p12113);
FA fa3870(ip_60_61,ip_61_60,ip_62_59,p12114,p12115);
FA fa3871(ip_63_58,p12113,p12092,p12116,p12117);
HA ha2187(p12115,p12088,p12118,p12119);
FA fa3872(p12090,p12094,p12117,p12120,p12121);
HA ha2188(p12096,p12098,p12122,p12123);
HA ha2189(p12119,p12100,p12124,p12125);
FA fa3873(p12121,p12123,p12125,p12126,p12127);
FA fa3874(p12127,p12102,p12104,p12128,p12129);
FA fa3875(p12106,p12108,p12129,p12130,p12131);
HA ha2190(ip_59_63,ip_60_62,p12132,p12133);
HA ha2191(ip_61_61,ip_62_60,p12134,p12135);
HA ha2192(ip_63_59,p12112,p12136,p12137);
HA ha2193(p12133,p12135,p12138,p12139);
HA ha2194(p12137,p12139,p12140,p12141);
HA ha2195(p12114,p12141,p12142,p12143);
FA fa3876(p12116,p12118,p12143,p12144,p12145);
FA fa3877(p12122,p12120,p12124,p12146,p12147);
HA ha2196(p12145,p12126,p12148,p12149);
FA fa3878(p12147,p12149,p12128,p12150,p12151);
HA ha2197(ip_60_63,ip_61_62,p12152,p12153);
HA ha2198(ip_62_61,ip_63_60,p12154,p12155);
HA ha2199(p12132,p12134,p12156,p12157);
FA fa3879(p12153,p12155,p12136,p12158,p12159);
HA ha2200(p12138,p12157,p12160,p12161);
HA ha2201(p12140,p12159,p12162,p12163);
HA ha2202(p12161,p12142,p12164,p12165);
FA fa3880(p12163,p12165,p12144,p12166,p12167);
FA fa3881(p12167,p12146,p12148,p12168,p12169);
FA fa3882(ip_61_63,ip_62_62,ip_63_61,p12170,p12171);
FA fa3883(p12152,p12154,p12156,p12172,p12173);
FA fa3884(p12171,p12160,p12173,p12174,p12175);
FA fa3885(p12158,p12162,p12164,p12176,p12177);
HA ha2203(p12175,p12177,p12178,p12179);
HA ha2204(p12179,p12166,p12180,p12181);
FA fa3886(ip_62_63,ip_63_62,p12170,p12182,p12183);
HA ha2205(p12172,p12183,p12184,p12185);
FA fa3887(p12185,p12174,p12176,p12186,p12187);
HA ha2206(p12178,p12187,p12188,p12189);
FA fa3888(ip_63_63,p12182,p12184,p12190,p12191);
HA ha2207(p12191,p12186,p12192,p12193);
wire [127:0] a,b;
wire [127:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = ip_2_0;
assign b[2] = p1;
assign a[3] = p5;
assign b[3] = 1'b0;
assign a[4] = p11;
assign b[4] = 1'b0;
assign a[5] = p19;
assign b[5] = 1'b0;
assign a[6] = p31;
assign b[6] = 1'b0;
assign a[7] = p43;
assign b[7] = p30;
assign a[8] = p59;
assign b[8] = 1'b0;
assign a[9] = p77;
assign b[9] = 1'b0;
assign a[10] = p103;
assign b[10] = p76;
assign a[11] = p102;
assign b[11] = p131;
assign a[12] = p163;
assign b[12] = p130;
assign a[13] = p193;
assign b[13] = p195;
assign a[14] = p233;
assign b[14] = p194;
assign a[15] = p275;
assign b[15] = p232;
assign a[16] = p315;
assign b[16] = 1'b0;
assign a[17] = p359;
assign b[17] = p314;
assign a[18] = p407;
assign b[18] = 1'b0;
assign a[19] = p463;
assign b[19] = p406;
assign a[20] = p517;
assign b[20] = 1'b0;
assign a[21] = p575;
assign b[21] = p516;
assign a[22] = p637;
assign b[22] = 1'b0;
assign a[23] = p701;
assign b[23] = 1'b0;
assign a[24] = p773;
assign b[24] = p700;
assign a[25] = p772;
assign b[25] = p845;
assign a[26] = p913;
assign b[26] = p844;
assign a[27] = p991;
assign b[27] = 1'b0;
assign a[28] = p1065;
assign b[28] = p990;
assign a[29] = p1149;
assign b[29] = 1'b0;
assign a[30] = p1229;
assign b[30] = p1148;
assign a[31] = p1321;
assign b[31] = 1'b0;
assign a[32] = p1411;
assign b[32] = 1'b0;
assign a[33] = p1505;
assign b[33] = p1410;
assign a[34] = p1504;
assign b[34] = p1603;
assign a[35] = p1705;
assign b[35] = p1602;
assign a[36] = p1704;
assign b[36] = p1809;
assign a[37] = p1911;
assign b[37] = p1808;
assign a[38] = p2017;
assign b[38] = 1'b0;
assign a[39] = p2125;
assign b[39] = p2016;
assign a[40] = p2241;
assign b[40] = 1'b0;
assign a[41] = p2363;
assign b[41] = p2240;
assign a[42] = p2491;
assign b[42] = 1'b0;
assign a[43] = p2619;
assign b[43] = p2490;
assign a[44] = p2618;
assign b[44] = p2753;
assign a[45] = p2897;
assign b[45] = 1'b0;
assign a[46] = p3037;
assign b[46] = p2896;
assign a[47] = p3175;
assign b[47] = 1'b0;
assign a[48] = p3323;
assign b[48] = p3174;
assign a[49] = p3322;
assign b[49] = p3473;
assign a[50] = p3472;
assign b[50] = p3623;
assign a[51] = p3771;
assign b[51] = p3622;
assign a[52] = p3770;
assign b[52] = p3919;
assign a[53] = p4065;
assign b[53] = p3918;
assign a[54] = p4064;
assign b[54] = p4221;
assign a[55] = p4381;
assign b[55] = 1'b0;
assign a[56] = p4547;
assign b[56] = p4380;
assign a[57] = p4546;
assign b[57] = p4721;
assign a[58] = p4901;
assign b[58] = p4720;
assign a[59] = p5089;
assign b[59] = 1'b0;
assign a[60] = p5289;
assign b[60] = p5088;
assign a[61] = p5288;
assign b[61] = p5487;
assign a[62] = p5689;
assign b[62] = 1'b0;
assign a[63] = p5881;
assign b[63] = p5688;
assign a[64] = p6073;
assign b[64] = 1'b0;
assign a[65] = p6257;
assign b[65] = 1'b0;
assign a[66] = p6441;
assign b[66] = 1'b0;
assign a[67] = p6623;
assign b[67] = p6440;
assign a[68] = p6807;
assign b[68] = 1'b0;
assign a[69] = p6977;
assign b[69] = p6806;
assign a[70] = p7145;
assign b[70] = p6976;
assign a[71] = p7319;
assign b[71] = 1'b0;
assign a[72] = p7491;
assign b[72] = p7318;
assign a[73] = p7665;
assign b[73] = 1'b0;
assign a[74] = p7835;
assign b[74] = 1'b0;
assign a[75] = p7991;
assign b[75] = p7834;
assign a[76] = p8149;
assign b[76] = 1'b0;
assign a[77] = p8303;
assign b[77] = 1'b0;
assign a[78] = p8457;
assign b[78] = 1'b0;
assign a[79] = p8609;
assign b[79] = 1'b0;
assign a[80] = p8759;
assign b[80] = p8608;
assign a[81] = p8903;
assign b[81] = p8758;
assign a[82] = p9039;
assign b[82] = 1'b0;
assign a[83] = p9169;
assign b[83] = 1'b0;
assign a[84] = p9303;
assign b[84] = 1'b0;
assign a[85] = p9431;
assign b[85] = 1'b0;
assign a[86] = p9557;
assign b[86] = 1'b0;
assign a[87] = p9691;
assign b[87] = p9556;
assign a[88] = p9819;
assign b[88] = p9690;
assign a[89] = p9937;
assign b[89] = 1'b0;
assign a[90] = p10057;
assign b[90] = 1'b0;
assign a[91] = p10165;
assign b[91] = p10056;
assign a[92] = p10281;
assign b[92] = p10164;
assign a[93] = p10391;
assign b[93] = 1'b0;
assign a[94] = p10495;
assign b[94] = p10390;
assign a[95] = p10601;
assign b[95] = p10494;
assign a[96] = p10600;
assign b[96] = p10701;
assign a[97] = p10805;
assign b[97] = p10700;
assign a[98] = p10804;
assign b[98] = p10901;
assign a[99] = p10900;
assign b[99] = p10993;
assign a[100] = p11077;
assign b[100] = 1'b0;
assign a[101] = p11157;
assign b[101] = p11076;
assign a[102] = p11239;
assign b[102] = 1'b0;
assign a[103] = p11319;
assign b[103] = p11238;
assign a[104] = p11389;
assign b[104] = p11318;
assign a[105] = p11388;
assign b[105] = p11457;
assign a[106] = p11456;
assign b[106] = p11521;
assign a[107] = p11587;
assign b[107] = 1'b0;
assign a[108] = p11649;
assign b[108] = 1'b0;
assign a[109] = p11703;
assign b[109] = p11648;
assign a[110] = p11763;
assign b[110] = 1'b0;
assign a[111] = p11815;
assign b[111] = p11762;
assign a[112] = p11861;
assign b[112] = p11814;
assign a[113] = p11903;
assign b[113] = p11860;
assign a[114] = p11902;
assign b[114] = p11939;
assign a[115] = p11973;
assign b[115] = 1'b0;
assign a[116] = p12003;
assign b[116] = p11972;
assign a[117] = p12033;
assign b[117] = p12002;
assign a[118] = p12061;
assign b[118] = p12032;
assign a[119] = p12087;
assign b[119] = p12060;
assign a[120] = p12086;
assign b[120] = p12111;
assign a[121] = p12131;
assign b[121] = p12110;
assign a[122] = p12151;
assign b[122] = p12130;
assign a[123] = p12169;
assign b[123] = p12150;
assign a[124] = p12181;
assign b[124] = p12168;
assign a[125] = p12189;
assign b[125] = p12180;
assign a[126] = p12188;
assign b[126] = p12193;
assign a[127] = p12190;
assign b[127] = p12192;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[127] = s[127];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
assign o[15] = s[15];
assign o[16] = s[16];
assign o[17] = s[17];
assign o[18] = s[18];
assign o[19] = s[19];
assign o[20] = s[20];
assign o[21] = s[21];
assign o[22] = s[22];
assign o[23] = s[23];
assign o[24] = s[24];
assign o[25] = s[25];
assign o[26] = s[26];
assign o[27] = s[27];
assign o[28] = s[28];
assign o[29] = s[29];
assign o[30] = s[30];
assign o[31] = s[31];
assign o[32] = s[32];
assign o[33] = s[33];
assign o[34] = s[34];
assign o[35] = s[35];
assign o[36] = s[36];
assign o[37] = s[37];
assign o[38] = s[38];
assign o[39] = s[39];
assign o[40] = s[40];
assign o[41] = s[41];
assign o[42] = s[42];
assign o[43] = s[43];
assign o[44] = s[44];
assign o[45] = s[45];
assign o[46] = s[46];
assign o[47] = s[47];
assign o[48] = s[48];
assign o[49] = s[49];
assign o[50] = s[50];
assign o[51] = s[51];
assign o[52] = s[52];
assign o[53] = s[53];
assign o[54] = s[54];
assign o[55] = s[55];
assign o[56] = s[56];
assign o[57] = s[57];
assign o[58] = s[58];
assign o[59] = s[59];
assign o[60] = s[60];
assign o[61] = s[61];
assign o[62] = s[62];
assign o[63] = s[63];
assign o[64] = s[64];
assign o[65] = s[65];
assign o[66] = s[66];
assign o[67] = s[67];
assign o[68] = s[68];
assign o[69] = s[69];
assign o[70] = s[70];
assign o[71] = s[71];
assign o[72] = s[72];
assign o[73] = s[73];
assign o[74] = s[74];
assign o[75] = s[75];
assign o[76] = s[76];
assign o[77] = s[77];
assign o[78] = s[78];
assign o[79] = s[79];
assign o[80] = s[80];
assign o[81] = s[81];
assign o[82] = s[82];
assign o[83] = s[83];
assign o[84] = s[84];
assign o[85] = s[85];
assign o[86] = s[86];
assign o[87] = s[87];
assign o[88] = s[88];
assign o[89] = s[89];
assign o[90] = s[90];
assign o[91] = s[91];
assign o[92] = s[92];
assign o[93] = s[93];
assign o[94] = s[94];
assign o[95] = s[95];
assign o[96] = s[96];
assign o[97] = s[97];
assign o[98] = s[98];
assign o[99] = s[99];
assign o[100] = s[100];
assign o[101] = s[101];
assign o[102] = s[102];
assign o[103] = s[103];
assign o[104] = s[104];
assign o[105] = s[105];
assign o[106] = s[106];
assign o[107] = s[107];
assign o[108] = s[108];
assign o[109] = s[109];
assign o[110] = s[110];
assign o[111] = s[111];
assign o[112] = s[112];
assign o[113] = s[113];
assign o[114] = s[114];
assign o[115] = s[115];
assign o[116] = s[116];
assign o[117] = s[117];
assign o[118] = s[118];
assign o[119] = s[119];
assign o[120] = s[120];
assign o[121] = s[121];
assign o[122] = s[122];
assign o[123] = s[123];
assign o[124] = s[124];
assign o[125] = s[125];
assign o[126] = s[126];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [127:0] a,b;
output [127:0] s;
assign s = a+b;
endmodule
