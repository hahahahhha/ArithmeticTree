// 1 2 1 2 2 1 2 2 2 1 2 1 2 1 1 2 

module main(x,y,o);
input [7:0] x,y;
output [15:0] o;
wire ip_0_0,ip_0_1,ip_0_2,ip_0_3,ip_0_4,ip_0_5,ip_0_6,ip_0_7,ip_1_0,ip_1_1,ip_1_2,ip_1_3,ip_1_4,ip_1_5,ip_1_6,ip_1_7,ip_2_0,ip_2_1,ip_2_2,ip_2_3,ip_2_4,ip_2_5,ip_2_6,ip_2_7,ip_3_0,ip_3_1,ip_3_2,ip_3_3,ip_3_4,ip_3_5,ip_3_6,ip_3_7,ip_4_0,ip_4_1,ip_4_2,ip_4_3,ip_4_4,ip_4_5,ip_4_6,ip_4_7,ip_5_0,ip_5_1,ip_5_2,ip_5_3,ip_5_4,ip_5_5,ip_5_6,ip_5_7,ip_6_0,ip_6_1,ip_6_2,ip_6_3,ip_6_4,ip_6_5,ip_6_6,ip_6_7,ip_7_0,ip_7_1,ip_7_2,ip_7_3,ip_7_4,ip_7_5,ip_7_6,ip_7_7;
wire p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63,p64,p65,p66,p67,p68,p69,p70,p71,p72,p73,p74,p75,p76,p77,p78,p79,p80,p81,p82,p83,p84,p85,p86,p87,p88,p89,p90,p91,p92,p93,p94,p95,p96,p97,p98,p99,p100,p101,p102,p103,p104,p105,p106,p107,p108,p109,p110,p111,p112,p113,p114,p115,p116,p117;
and and0(ip_0_0,x[0],y[0]);
and and1(ip_0_1,x[0],y[1]);
and and2(ip_0_2,x[0],y[2]);
and and3(ip_0_3,x[0],y[3]);
and and4(ip_0_4,x[0],y[4]);
and and5(ip_0_5,x[0],y[5]);
and and6(ip_0_6,x[0],y[6]);
and and7(ip_0_7,x[0],y[7]);
and and8(ip_1_0,x[1],y[0]);
and and9(ip_1_1,x[1],y[1]);
and and10(ip_1_2,x[1],y[2]);
and and11(ip_1_3,x[1],y[3]);
and and12(ip_1_4,x[1],y[4]);
and and13(ip_1_5,x[1],y[5]);
and and14(ip_1_6,x[1],y[6]);
and and15(ip_1_7,x[1],y[7]);
and and16(ip_2_0,x[2],y[0]);
and and17(ip_2_1,x[2],y[1]);
and and18(ip_2_2,x[2],y[2]);
and and19(ip_2_3,x[2],y[3]);
and and20(ip_2_4,x[2],y[4]);
and and21(ip_2_5,x[2],y[5]);
and and22(ip_2_6,x[2],y[6]);
and and23(ip_2_7,x[2],y[7]);
and and24(ip_3_0,x[3],y[0]);
and and25(ip_3_1,x[3],y[1]);
and and26(ip_3_2,x[3],y[2]);
and and27(ip_3_3,x[3],y[3]);
and and28(ip_3_4,x[3],y[4]);
and and29(ip_3_5,x[3],y[5]);
and and30(ip_3_6,x[3],y[6]);
and and31(ip_3_7,x[3],y[7]);
and and32(ip_4_0,x[4],y[0]);
and and33(ip_4_1,x[4],y[1]);
and and34(ip_4_2,x[4],y[2]);
and and35(ip_4_3,x[4],y[3]);
and and36(ip_4_4,x[4],y[4]);
and and37(ip_4_5,x[4],y[5]);
and and38(ip_4_6,x[4],y[6]);
and and39(ip_4_7,x[4],y[7]);
and and40(ip_5_0,x[5],y[0]);
and and41(ip_5_1,x[5],y[1]);
and and42(ip_5_2,x[5],y[2]);
and and43(ip_5_3,x[5],y[3]);
and and44(ip_5_4,x[5],y[4]);
and and45(ip_5_5,x[5],y[5]);
and and46(ip_5_6,x[5],y[6]);
and and47(ip_5_7,x[5],y[7]);
and and48(ip_6_0,x[6],y[0]);
and and49(ip_6_1,x[6],y[1]);
and and50(ip_6_2,x[6],y[2]);
and and51(ip_6_3,x[6],y[3]);
and and52(ip_6_4,x[6],y[4]);
and and53(ip_6_5,x[6],y[5]);
and and54(ip_6_6,x[6],y[6]);
and and55(ip_6_7,x[6],y[7]);
and and56(ip_7_0,x[7],y[0]);
and and57(ip_7_1,x[7],y[1]);
and and58(ip_7_2,x[7],y[2]);
and and59(ip_7_3,x[7],y[3]);
and and60(ip_7_4,x[7],y[4]);
and and61(ip_7_5,x[7],y[5]);
and and62(ip_7_6,x[7],y[6]);
and and63(ip_7_7,x[7],y[7]);
FA fa0(ip_0_2,ip_1_1,ip_2_0,p0,p1);
FA fa1(ip_0_3,ip_1_2,ip_2_1,p2,p3);
HA ha0(ip_3_0,p3,p4,p5);
FA fa2(ip_0_4,ip_1_3,ip_2_2,p6,p7);
HA ha1(ip_3_1,ip_4_0,p8,p9);
FA fa3(p9,p7,p2,p10,p11);
FA fa4(ip_0_5,ip_1_4,ip_2_3,p12,p13);
HA ha2(ip_3_2,ip_4_1,p14,p15);
FA fa5(ip_5_0,p15,p8,p16,p17);
HA ha3(p13,p17,p18,p19);
FA fa6(p6,p19,p10,p20,p21);
FA fa7(ip_0_6,ip_1_5,ip_2_4,p22,p23);
FA fa8(ip_3_3,ip_4_2,ip_5_1,p24,p25);
FA fa9(ip_6_0,p14,p23,p26,p27);
FA fa10(p25,p12,p27,p28,p29);
FA fa11(p16,p18,p29,p30,p31);
FA fa12(ip_0_7,ip_1_6,ip_2_5,p32,p33);
HA ha4(ip_3_4,ip_4_3,p34,p35);
FA fa13(ip_5_2,ip_6_1,ip_7_0,p36,p37);
FA fa14(p35,p33,p37,p38,p39);
FA fa15(p22,p24,p26,p40,p41);
FA fa16(p39,p41,p28,p42,p43);
HA ha5(ip_1_7,ip_2_6,p44,p45);
FA fa17(ip_3_5,ip_4_4,ip_5_3,p46,p47);
HA ha6(ip_6_2,ip_7_1,p48,p49);
FA fa18(p34,p45,p49,p50,p51);
HA ha7(p47,p32,p52,p53);
FA fa19(p36,p51,p53,p54,p55);
FA fa20(p38,p55,p40,p56,p57);
FA fa21(ip_2_7,ip_3_6,ip_4_5,p58,p59);
FA fa22(ip_5_4,ip_6_3,ip_7_2,p60,p61);
HA ha8(p44,p48,p62,p63);
FA fa23(p59,p61,p63,p64,p65);
HA ha9(p46,p50,p66,p67);
FA fa24(p52,p65,p67,p68,p69);
FA fa25(p54,p69,p56,p70,p71);
FA fa26(ip_3_7,ip_4_6,ip_5_5,p72,p73);
HA ha10(ip_6_4,ip_7_3,p74,p75);
HA ha11(p75,p62,p76,p77);
FA fa27(p73,p58,p60,p78,p79);
HA ha12(p77,p64,p80,p81);
HA ha13(p66,p79,p82,p83);
FA fa28(p81,p83,p68,p84,p85);
FA fa29(ip_4_7,ip_5_6,ip_6_5,p86,p87);
FA fa30(ip_7_4,p74,p87,p88,p89);
FA fa31(p72,p76,p89,p90,p91);
HA ha14(p91,p78,p92,p93);
HA ha15(p80,p82,p94,p95);
FA fa32(p93,p95,p84,p96,p97);
FA fa33(ip_5_7,ip_6_6,ip_7_5,p98,p99);
HA ha16(p99,p86,p100,p101);
FA fa34(p101,p88,p90,p102,p103);
HA ha17(p103,p92,p104,p105);
HA ha18(p94,p105,p106,p107);
FA fa35(ip_6_7,ip_7_6,p98,p108,p109);
FA fa36(p100,p109,p102,p110,p111);
FA fa37(p104,p106,p111,p112,p113);
HA ha19(ip_7_7,p108,p114,p115);
FA fa38(p115,p110,p112,p116,p117);
wire [15:0] a,b;
wire [15:0] s;
assign a[1] = ip_0_1;
assign b[1] = ip_1_0;
assign a[2] = p1;
assign b[2] = 1'b0;
assign a[3] = p0;
assign b[3] = p5;
assign a[4] = p4;
assign b[4] = p11;
assign a[5] = p21;
assign b[5] = 1'b0;
assign a[6] = p31;
assign b[6] = p20;
assign a[7] = p30;
assign b[7] = p43;
assign a[8] = p57;
assign b[8] = p42;
assign a[9] = p71;
assign b[9] = 1'b0;
assign a[10] = p85;
assign b[10] = p70;
assign a[11] = p97;
assign b[11] = 1'b0;
assign a[12] = p107;
assign b[12] = p96;
assign a[13] = p113;
assign b[13] = 1'b0;
assign a[14] = p117;
assign b[14] = 1'b0;
assign a[15] = p114;
assign b[15] = p116;
assign a[0] = ip_0_0;
assign b[0] = 1'b0;
assign o[15] = s[15];
assign o[0] = s[0];
assign o[1] = s[1];
assign o[2] = s[2];
assign o[3] = s[3];
assign o[4] = s[4];
assign o[5] = s[5];
assign o[6] = s[6];
assign o[7] = s[7];
assign o[8] = s[8];
assign o[9] = s[9];
assign o[10] = s[10];
assign o[11] = s[11];
assign o[12] = s[12];
assign o[13] = s[13];
assign o[14] = s[14];
adder add(a,b,s);

endmodule

module HA(a,b,c,s);
input a,b;
output c,s;
xor x1(s,a,b);
and a1(c,a,b);
endmodule
module FA(a,b,c,cy,sm);
input a,b,c;
output cy,sm;
wire x,y,z;
HA h1(a,b,x,z);
HA h2(z,c,y,sm);
or o1(cy,x,y);
endmodule

module adder(a,b,s);
input [15:0] a,b;
output [15:0] s;
assign s = a+b;
endmodule
